-- File:        OrientedFace.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWOrientedFace from RWStepShape

	---Purpose : Read & Write Module for OrientedFace

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     OrientedFace from StepShape,
     EntityIterator from Interface

is

	Create returns RWOrientedFace;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable OrientedFace from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : OrientedFace from StepShape);

	Share(me; ent : OrientedFace from StepShape; iter : in out EntityIterator);

end RWOrientedFace;
