-- File:        RectangularCompositeSurface.cdl
-- Created:     Mon Dec  4 12:02:30 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWRectangularCompositeSurface from RWStepGeom

	---Purpose : Read & Write Module for RectangularCompositeSurface

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     RectangularCompositeSurface from StepGeom,
     EntityIterator from Interface

is

	Create returns RWRectangularCompositeSurface;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable RectangularCompositeSurface from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : RectangularCompositeSurface from StepGeom);

	Share(me; ent : RectangularCompositeSurface from StepGeom; iter : in out EntityIterator);

end RWRectangularCompositeSurface;
