-- File:	RWStepFEA_RWFeaMoistureAbsorption.cdl
-- Created:	Thu Dec 12 17:51:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFeaMoistureAbsorption from RWStepFEA

    ---Purpose: Read & Write tool for FeaMoistureAbsorption

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FeaMoistureAbsorption from StepFEA

is
    Create returns RWFeaMoistureAbsorption from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FeaMoistureAbsorption from StepFEA);
	---Purpose: Reads FeaMoistureAbsorption

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FeaMoistureAbsorption from StepFEA);
	---Purpose: Writes FeaMoistureAbsorption

    Share (me; ent : FeaMoistureAbsorption from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFeaMoistureAbsorption;
