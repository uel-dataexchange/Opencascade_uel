-- File:	Geom2d.cdl
-- Created:	Wed Mar 24 17:29:38 1993
-- Author:	JCV
--		<fid@sdsun2>
-- Copyright:	 Matra Datavision 1993

---Copyright:   Matra Datavision 1991


package Geom2d

        --- Purpose :
        --  This package contains the definition of the geometric objects 
        --  such as point, vector, axis placement, curves and the
        --  description of the geometric transformations available 
        --  for these objects.
        --  All these entities are defined in 2D space.
        --  This package gives the possibility :
        --     . to create geometric objects,
        --     . to have information about them,
        --     . to modify these objects.
        --  This package uses the services of the package gp (Geometric
        --  processor) which describes non-persistent objects for algebraic
        --  calculus and basic analytic geometry. The purpose of this package
        --  is to create persistent geometric objects and to read geometric
        --  information about these objects. Complexes geometric algorithmes
        --  are not described in this package.     At construction time,
        --  elementary verifications are done to verify that the objects
        --  are coherents, but some verifications which require complex
        --  algorithmes (for example to check that a curve has not null
        --  length or does not self-intersect) must be done before the 
        --  construction of the geometric objects. 


uses MMgt, GeomAbs, TColStd, gp, TColgp

is

exception UndefinedDerivative inherits DomainError  from  Standard;
exception UndefinedValue inherits DomainError   from  Standard ;



  class Transformation;


  deferred class Geometry;


     deferred class Point;
              class  CartesianPoint;


     deferred class Vector;
              class Direction;
              class VectorWithMagnitude;
     

     class AxisPlacement;


     deferred class Curve;

              class Line;

              deferred class Conic;
                       class Circle;
                       class Ellipse;
                       class Hyperbola;
                       class Parabola;

              deferred class BoundedCurve;
                       class BezierCurve;
                       class BSplineCurve;
                       class TrimmedCurve;

              class  OffsetCurve;


end Geom2d;




