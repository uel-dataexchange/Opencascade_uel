-- File:	PSurfaceTool.cdl
-- Created:	Fri Mar  6 16:32:01 1992
-- Author:	Isabelle GRIGNON
--		<isg@phobox>
---Copyright:	 Matra Datavision 1992


deferred generic class PSurfaceTool from IntImp
    (Surface as any)          
                                   

	---Purpose: Template class for a tool on a bi-parametrised surface.
	--          It is possible to implement this tool with an
	--          instantiation of the SurfaceTool from Adaptor3d.

uses Pnt from gp,
     Vec from gp
 
is

    UIntervalFirst(myclass ; S: Surface)
	   
	---Purpose: Returns the first U parameter of the surface.

    	returns Real from Standard;
    
    
    VIntervalFirst(myclass ; S: Surface)
	   
	---Purpose: Returns the first V parameter of the surface.

    	returns Real from Standard;
    
    
    UIntervalLast(myclass ; S: Surface)
	   
	---Purpose: Returns the last U parameter of the surface.

    	returns Real from Standard;
    
    
    VIntervalLast(myclass ; S: Surface)
	   
	---Purpose: Returns the last V parameter of the surface.

    	returns Real from Standard;
    
    
    Value (myclass ; S: Surface; U,V : Real from Standard)
    
    	---Purpose: Returns the point of parameter (U,V) on the surface.

    	returns Pnt from gp;


    D1(myclass; S: Surface; U,V: Real from Standard; 
                P: out Pnt from gp; D1U,D1V: out Vec from gp);
		
	---Purpose: Returns the point of parameter (U,V) on the surface,
	--          and the first derivatives in the directions u and v.

    
    UResolution(myclass; S : Surface; Tol3d: Real from Standard)
    
	---Purpose: Returns the numerical resolution in the U direction,
	--          for a given resolution in 3d space.

    	returns Real from Standard;


    VResolution(myclass; S : Surface; Tol3d: Real from Standard)
    
	---Purpose: Returns the numerical resolution in the V direction,
	--          for a given resolution in 3d space.

    	returns Real from Standard;


end PSurfaceTool;
