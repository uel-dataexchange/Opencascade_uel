-- File:        BoundedSurface.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWBoundedSurface from RWStepGeom

	---Purpose : Read & Write Module for BoundedSurface

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     BoundedSurface from StepGeom

is

	Create returns RWBoundedSurface;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable BoundedSurface from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : BoundedSurface from StepGeom);

end RWBoundedSurface;
