-- File:	RWStepDimTol_RWParallelismTolerance.cdl
-- Created:	Wed Jun  4 13:34:34 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWParallelismTolerance from RWStepDimTol

    ---Purpose: Read & Write tool for ParallelismTolerance

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ParallelismTolerance from StepDimTol

is
    Create returns RWParallelismTolerance from RWStepDimTol;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ParallelismTolerance from StepDimTol);
	---Purpose: Reads ParallelismTolerance

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ParallelismTolerance from StepDimTol);
	---Purpose: Writes ParallelismTolerance

    Share (me; ent : ParallelismTolerance from StepDimTol;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWParallelismTolerance;
