-- File:	IGESSolid_ToolVertexList.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolVertexList  from IGESSolid

    ---Purpose : Tool to work on a VertexList. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses VertexList from IGESSolid,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolVertexList;
    ---Purpose : Returns a ToolVertexList, ready to work


    ReadOwnParams (me; ent : mutable VertexList;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : VertexList;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : VertexList;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a VertexList <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : VertexList) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : VertexList;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : VertexList; entto : mutable VertexList;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : VertexList;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolVertexList;
