-- File:	RWStepRepr_RWSpecifiedHigherUsageOccurrence.cdl
-- Created:	Mon Jul  3 20:13:37 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWSpecifiedHigherUsageOccurrence from RWStepRepr

    ---Purpose: Read & Write tool for SpecifiedHigherUsageOccurrence

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    SpecifiedHigherUsageOccurrence from StepRepr

is
    Create returns RWSpecifiedHigherUsageOccurrence from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : SpecifiedHigherUsageOccurrence from StepRepr);
	---Purpose: Reads SpecifiedHigherUsageOccurrence

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: SpecifiedHigherUsageOccurrence from StepRepr);
	---Purpose: Writes SpecifiedHigherUsageOccurrence

    Share (me; ent : SpecifiedHigherUsageOccurrence from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWSpecifiedHigherUsageOccurrence;
