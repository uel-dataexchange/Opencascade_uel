-- File:	ToolPolyhedron.cdl
-- Created:	Wed Sep 18 08:44:42 1991
-- Author:	Didier PIFFAULT
--		<dpf@sdsun1>
---Copyright:	 Matra Datavision 1991, 1992


generic class ToolPolyhedron from Intf (Polyhedron as any)

    ---Purpose: Describes the signature  of  a polyedral surface with  only
    --          triangular facets and the information  necessary to compute
    --          the interferences.


uses    XYZ from gp,
    	Pnt from gp,
    	Box from Bnd,
	HArray1OfBox from Bnd


raises  OutOfRange from Standard


is  Bounding       (myclass; thePolyh : Polyhedron)
    	    	    returns Box from Bnd;
    ---Purpose: Returns the bounding box of the ToolPolyhedron.

    ComponentsBounding
       	    	   (myclass; thePolyh : Polyhedron)
    	    	    returns HArray1OfBox from Bnd;
    ---Purpose: Returns the array of boxes. The box <n> corresponding 
    --          to the triangle <n>.


    DeflectionOverEstimation
		   (myclass; thePolyh : Polyhedron)
    	    	    returns Real from Standard;
    ---Purpose: Returns the tolerance of the polygon.


-- Structure needings :

    NbTriangles	   (myclass; thePolyh : Polyhedron) 
    	    	    returns Integer from Standard;
    ---Purpose: Returns the number of triangles in this polyedron.


    Triangle	   (myclass; thePolyh : Polyhedron;
		    Index     : in Integer from Standard;
		    P1,P2,P3  : out Integer from Standard)
		    raises OutOfRange from Standard;
    ---Purpose: Returns the indices  of  the 3 points of  the triangle of
    --          address Index in the ToolPolyhedron.


    Point	   (myclass; thePolyh : Polyhedron;
		    Index : in Integer)
		    returns Pnt from gp
		    raises OutOfRange from Standard;
    ---Purpose: Returns the point of index i in the polyedron.


    TriConnex	   (myclass; thePolyh : Polyhedron;
		    Triang	 : in Integer;
		    Pivot,Pedge	 : in Integer;
		    TriCon	 : out Integer;
		    OtherPedge	 : out Integer)
		    returns Integer
		    raises OutOfRange from Standard;
    ---Purpose: Returns  the  triangle <Tricon> connected  to  the triangle
    --          <Triang> by  the edge <Pivot><Pedge>.   The  third point of
    --          the connected triangle is returned in <OtherPedge> (Used to
    --          turn  around a vertex).   When the edge  <Pivot><Pedge>  is
    --          free  (no  connected triangle) <Tricon> is  null.   In this
    --          case the function returns the triangle on the free bound of
    --          the polyhedron connected to <Triang> by vertex <Pivot>.



end ToolPolyhedron;
