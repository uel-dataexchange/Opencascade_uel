-- File:	GraphTools_GraphIterator.cdl
-- Created:	Wed Mar  6 18:20:11 1991
-- Author:	Denis Pascal
--		<dp@topsn3>
---Copyright:	 Matra Datavision 1991, 1992


generic class GraphIterator from GraphTools (Graph  as any;
				             Vertex as any)
				  
-- template class GraphIterator from GraphTools (Graph  as any;
--                                                Vertex as any)

    	---Purpose: Template  class which defines   signatures  of  an
    	--          iterator  to  visit  each  vertex,   member of the
    	--          underlying graph.


raises NoMoreObject from Standard,
       NoSuchObject from Standard

is

    Create (G : Graph) returns GraphIterator;

    More (me) returns Boolean;
	---Purpose: Returns TRUE if there are other vertices.
        ---Level: Public
    
    Next (me : in out)
    	--- Purpose : Set the iterator to the next Vertex.
        ---Level: Public
    raises NoMoreObject from Standard;

    Value (me) returns Vertex
	--- Purpose: Returns the vertex value for the current position
	--  of the iterator
        ---Level: Public
    raises NoSuchObject from Standard;

end GraphIterator;



















