-- File:	RWStepBasic_RWCertification.cdl
-- Created:	Fri Nov 26 16:26:34 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWCertification from RWStepBasic

    ---Purpose: Read & Write tool for Certification

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    Certification from StepBasic

is
    Create returns RWCertification from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : Certification from StepBasic);
	---Purpose: Reads Certification

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: Certification from StepBasic);
	---Purpose: Writes Certification

    Share (me; ent : Certification from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWCertification;
