-- File:	RWStepShape_RWEdgeBasedWireframeModel.cdl
-- Created:	Fri Dec 28 16:02:01 2001 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWEdgeBasedWireframeModel from RWStepShape

    ---Purpose: Read & Write tool for EdgeBasedWireframeModel

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    EdgeBasedWireframeModel from StepShape

is
    Create returns RWEdgeBasedWireframeModel from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : EdgeBasedWireframeModel from StepShape);
	---Purpose: Reads EdgeBasedWireframeModel

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: EdgeBasedWireframeModel from StepShape);
	---Purpose: Writes EdgeBasedWireframeModel

    Share (me; ent : EdgeBasedWireframeModel from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWEdgeBasedWireframeModel;
