-- File:        OrientedPath.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWOrientedPath from RWStepShape

	---Purpose : Read & Write Module for OrientedPath

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     OrientedPath from StepShape,
     EntityIterator from Interface

is

	Create returns RWOrientedPath;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable OrientedPath from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : OrientedPath from StepShape);

	Share(me; ent : OrientedPath from StepShape; iter : in out EntityIterator);

end RWOrientedPath;
