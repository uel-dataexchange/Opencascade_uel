-- File:	RWStepAP214_RWExternallyDefinedClass.cdl
-- Created:	Wed May 10 15:09:06 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWExternallyDefinedClass from RWStepAP214

    ---Purpose: Read & Write tool for ExternallyDefinedClass

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ExternallyDefinedClass from StepAP214

is
    Create returns RWExternallyDefinedClass from RWStepAP214;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ExternallyDefinedClass from StepAP214);
	---Purpose: Reads ExternallyDefinedClass

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ExternallyDefinedClass from StepAP214);
	---Purpose: Writes ExternallyDefinedClass

    Share (me; ent : ExternallyDefinedClass from StepAP214;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWExternallyDefinedClass;
