-- File:	TDF_RelocationTable.cdl
--      	-----------------------
-- Author:	DAUTRY Philippe
--		<fid@fox.paris1.matra-dtv.fr>
---Copyright:	 MATRA DATAVISION 1997

---Version:	0.0
---History:	Version	Date		Purpose
--		0.0	Mar  6 1997	Creation
--		1.0	Sep 23 1998	DoubleMaps->DataMap


class RelocationTable from TDF
    inherits TShared from MMgt

	---Purpose: This is a relocation dictionnary between source
	--          and target labels, attributes or any
	--          transient. Note that one target value may be the
	--          relocation value of more than one source object.
	--          
	--          Common behaviour: it returns true and the found
	--          relocation value as target object; false
	--          otherwise.
	--          
	--          Look at SelfRelocate method for more explanation
	--          about self relocation behavior of this class.


uses

    Attribute           from TDF,
    Data                from TDF,
    Label               from TDF,
    LabelMap            from TDF,
    LabelDataMap        from TDF,
    AttributeMap        from TDF,
    AttributeDataMap    from TDF,
    IndexedDataMapOfTransientTransient from TColStd

-- raises

is

    Create(selfRelocate : Boolean from Standard = Standard_False)
--    Create(selfRelocate : Boolean from Standard = Standard_False;afterRelocate :Boolean from Standard = Standard_False)     
    	returns mutable RelocationTable from TDF;
	---Purpose: Creates an relocation table. <selfRelocate> says
	--          if a value without explicit relocation is its own
	--          relocation.


    ---Category: Self relocation methods.
    --           -------------------------

    SelfRelocate(me : mutable; selfRelocate : Boolean from Standard);
	---Purpose: Sets <mySelfRelocate> to <selfRelocate>.
	--          
	--          This flag affects the HasRelocation method
	--          behavior like this:
	--          
	--          <mySelfRelocate> == False:
	--          
	--          If no relocation object is found in the map, a
	--          null object is returned
	--          
	--          <mySelfRelocate> == True:
	--          
	--          If no relocation object is found in the map, the
	--          method assumes the source object is relocation
	--          value; so the source object is returned as target
	--          object.

    SelfRelocate(me) returns Boolean from Standard;
	---Purpose: Returns <mySelfRelocate>.

    AfterRelocate(me : mutable; afterRelocate : Boolean from Standard);

    AfterRelocate(me) returns Boolean from Standard;
	---Purpose: Returns <myAfterRelocate>.

    ---Category: Label relocation methods.
    --           -------------------------

    SetRelocation(me : mutable;
    	       	  aSourceLabel : Label from TDF;
    	       	  aTargetLabel : Label from TDF);
	---Purpose: Sets the relocation value of <aSourceLabel> to
	--          <aTargetLabel>.

    HasRelocation(me;
    	     	  aSourceLabel :        Label from TDF;
    	     	  aTargetLabel : in out Label from TDF)
	returns Boolean from Standard;
	---Purpose: Finds the relocation value of <aSourceLabel>
	--          and returns it into <aTargetLabel>.
	--          
	--          (See above SelfRelocate method for more
	--          explanation about the method behavior)


    ---Category: Attribute relocation methods.
    --           -----------------------------

    SetRelocation(me : mutable;
    	       	  aSourceAttribute : Attribute from TDF;
    	       	  aTargetAttribute : Attribute from TDF);
	---Purpose: Sets the relocation value of <aSourceAttribute> to
	--          <aTargetAttribute>.

    HasRelocation(me;
    	     	  aSourceAttribute :               Attribute from TDF;
    	     	  aTargetAttribute : in out mutable Attribute from TDF)
	returns Boolean from Standard;
	---Purpose: Finds the relocation value of <aSourceAttribute>
	--          and returns it into <aTargetAttribute>.
	--          
	--          (See above SelfRelocate method for more
	--          explanation about the method behavior)


    ---Category: Transient other types object relocation methods.
    --           ------------------------------------------------

    SetTransientRelocation(me : mutable;
    	                   aSourceTransient : Transient from Standard;
    	                   aTargetTransient : Transient from Standard);
	---Purpose: Sets the relocation value of <aSourceTransient> to
	--          <aTargetTransient>.

    HasTransientRelocation
    	(me;
    	 aSourceTransient :                Transient from Standard;
    	 aTargetTransient : in out mutable Transient from Standard)
	returns Boolean from Standard;
	---Purpose: Finds the relocation value of <aSourceTransient>
	--          and returns it into <aTargetTransient>.
	--          
	--          (See above SelfRelocate method for more
	--          explanation about the method behavior)

    ---Category: Miscelleaneous
    --           --------------

    Clear(me : mutable);
	---Purpose: Clears the relocation dictionnary, but lets the
	--          self relocation flag to its current value.

    TargetLabelMap(me; aLabelMap : in out LabelMap from TDF);
	---Purpose: Fills <aLabelMap> with target relocation
	--          labels. <aLabelMap> is not cleared before use.

    TargetAttributeMap(me; anAttributeMap : in out AttributeMap from TDF);
	---Purpose: Fills <anAttributeMap> with target relocation
	--          attributes. <anAttributeMap> is not cleared before
	--          use.

    -- Try not to use the following methods, for they are very
    -- implementation dependent.

    LabelTable(me : mutable)
    	returns LabelDataMap from TDF;
	---Purpose: Returns <myLabelTable> to be used or updated.
	--          
	---C++: return &

    AttributeTable(me : mutable)
    	returns AttributeDataMap from TDF;
	---Purpose: Returns <myAttributeTable> to be used or updated.
	--          
	---C++: return &

    TransientTable(me : mutable)
    	returns IndexedDataMapOfTransientTransient from TColStd;
	---Purpose: Returns <myTransientTable> to be used or updated.
	--          
	---C++: return &

    Dump(me;
    	 dumpLabels, dumpAttributes, dumpTransients : Boolean from Standard;
	 anOS : in out OStream from Standard)
    	returns OStream from Standard;
	---Purpose: Dumps the relocation table.
	--          
	---C++: return &

fields

    mySelfRelocate    : Boolean from Standard;
    myAfterRelocate   : Boolean from Standard;
    myLabelTable      : LabelDataMap     from TDF;
    myAttributeTable  : AttributeDataMap from TDF;
    myTransientTable  : IndexedDataMapOfTransientTransient from TColStd;
    -- Indexed... because there is no other type available in TColStd.

end RelocationTable from TDF;
