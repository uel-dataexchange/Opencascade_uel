-- File:        BinMDataStd_RealListDriver.cdl
-- Created:     May 29 11:40:00 2007
-- Author:      Vlad Romashko
--  	    	<vladislav.romashko@opencascade.com>
-- Copyright:   Open CASCADE

class RealListDriver from BinMDataStd inherits ADriver from BinMDF

uses

    MessageDriver    from CDM,
    SRelocationTable from BinObjMgt,
    RRelocationTable from BinObjMgt,
    Persistent       from BinObjMgt,
    Attribute        from TDF

is
    Create (theMessageDriver:MessageDriver from CDM)
    returns mutable RealListDriver from BinMDataStd;

    NewEmpty (me)
    returns mutable Attribute from TDF
    is redefined;

    Paste(me; Source     : Persistent from BinObjMgt;
              Target     : mutable Attribute from TDF;
              RelocTable : out RRelocationTable from BinObjMgt)
    returns Boolean from Standard is redefined;

    Paste(me; Source     : Attribute from TDF;
              Target     : in out Persistent from BinObjMgt;
              RelocTable : out SRelocationTable from BinObjMgt)
    is redefined;

end RealListDriver;
