-- File:        RightAngularWedge.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWRightAngularWedge from RWStepShape

	---Purpose : Read & Write Module for RightAngularWedge

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     RightAngularWedge from StepShape,
     EntityIterator from Interface

is

	Create returns RWRightAngularWedge;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable RightAngularWedge from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : RightAngularWedge from StepShape);

	Share(me; ent : RightAngularWedge from StepShape; iter : in out EntityIterator);

end RWRightAngularWedge;
