-- File:	GeomFill_SnglrFunc.cdl
-- Created:	Thu Feb 26 10:42:27 1998
-- Author:	Roman BORISOV
--		<rbv@ecolox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1998


private class SnglrFunc from GeomFill inherits  Curve  from  Adaptor3d

	---Purpose: to  represent  function  C'(t)^C''(t)

uses
    HCurve from Adaptor3d, 
    Shape  from GeomAbs, 
    CurveType  from GeomAbs,
    Array1OfReal from TColStd, 
    Pnt from gp, 
    Vec from gp
    
raises
    OutOfRange from Standard, 
    DomainError from Standard

is
    Create(HC: HCurve from Adaptor3d) 
      returns SnglrFunc;  
       
    SetRatio(me:in  out;  Ratio  :  Real) 
      is  static;
   
    FirstParameter(me) returns Real
      is redefined static;

    LastParameter(me) returns Real
      is redefined static; 
     
    NbIntervals(me: in out; S : Shape from GeomAbs) returns Integer
	---Purpose: Returns  the number  of  intervals for  continuity
	--          <S>. May be one if Continuity(me) >= <S>
    is redefined static;
    
    Intervals(me: in out; T : in out Array1OfReal from TColStd; 
    	          S : Shape from GeomAbs)
	---Purpose: Stores in <T> the  parameters bounding the intervals
	--          of continuity <S>.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
    raises
    	OutOfRange from Standard 
    is redefined static;  

    Value(me; U : Real) returns Pnt from gp
         --- Purpose : Computes the point of parameter U on the curve.
    is redefined static;
 
    IsPeriodic(me) returns Boolean
    is redefined static;
    
    Period(me) returns Real
    raises
    	DomainError from Standard -- if the curve is not periodic
    is redefined static;
    
    D0 (me; U : Real; P : out Pnt from gp)
         --- Purpose : Computes the point of parameter U on the curve.
    is redefined static;
    
    D1 (me; U : Real; P : out Pnt from gp ; V : out Vec from gp)
         --- Purpose : Computes the point of parameter U on the curve with its
         --  first derivative.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C1.
    is redefined static;
    
    D2 (me; U : Real; P : out Pnt from gp; V1, V2 : out Vec from gp)
        --- Purpose :
        --  Returns the point P of parameter U, the first and second
        --  derivatives V1 and V2.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C2.
     is redefined static;
 
    Resolution(me; R3d : Real) returns Real
         ---Purpose :  Returns the parametric  resolution corresponding
         --         to the real space resolution <R3d>.
    is redefined static;   

    GetType(me) returns CurveType from GeomAbs
	---Purpose: Returns  the  type of the   curve  in the  current
	--          interval :   Line,   Circle,   Ellipse, Hyperbola,
	--          Parabola, BezierCurve, BSplineCurve, OtherCurve.
    is redefined static;

fields 

  myHCurve: HCurve  from  Adaptor3d;  
  ratio   :  Real;
  
end SnglrFunc;
