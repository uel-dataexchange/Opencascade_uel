-- File:	Builder.cdl
-- Created:	Thu Mar 12 11:04:50 1992
-- Author:	Philippe DAUTRY
--		<fid@sdsun1>
---Copyright:	 Matra Datavision 1992



deferred generic class Builder from Primitives(
    TheShell  as any;
    TheFace   as any;
    TheWire   as any;
    TheEdge   as any;
    TheVertex as any)

	---Purpose: This is a signature class describing services from
	--          the  Topology Data   Structure   required  by  the
	--          Primitives algorithms.

uses
    Pnt      from gp,
    Lin      from gp,
    Circ     from gp,
    Pln      from gp,
    
    Lin2d    from gp,
    Circ2d   from gp

is
    MakeShell (me; S : out TheShell)
	---Purpose: Make a empty Shell.
    is deferred;
    
    MakeFace (me; F : out TheFace; P : Pln from gp)
	---Purpose: Returns in   <F> a  Face  built  with   the  plane
	--          equation <P>.
    is deferred;
    
    MakeWire(me; W : out TheWire)
	---Purpose: Returns in <W> an empty Wire.
    is deferred;
    
    MakeDegeneratedEdge (me; E : out TheEdge)
	---Purpose: Returns in <E> a degenerated edge.
    is deferred;

    MakeEdge (me; E : out TheEdge; L : Lin from gp)
	---Purpose: Returns   in <E>  an  Edge  built  with  the  line
	--          equation  <L>.
    is deferred;

    MakeEdge (me; E : out TheEdge; C : Circ from gp)
	---Purpose: Returns  in <E>   an  Edge  built  with the circle
	--          equation  <C>.
    is deferred;
    
    SetPCurve(me; E : in out TheEdge; F : in TheFace; L : Lin2d from gp)
	---Purpose: Sets the line <L> to be the curve representing the
	--          edge <E> in the parametric space of the surface of
	--          <F>.
    is deferred;
    
    SetPCurve(me; E : in out TheEdge; F : in TheFace; L1,L2 : Lin2d from gp)
	---Purpose: Sets the    lines  <L1,L2>  to   be     the curves
	--          representing the edge <E>  in the parametric space
	--          of the surface of <F>. The surface is closed.
    is deferred;
    
    SetPCurve(me; E : in out TheEdge; F : in TheFace; C : Circ2d from gp)
	---Purpose: Sets the  circle <C> to  be the curve representing
	--          the  edge <E>  in   the  parametric  space of  the
	--          surface of <F>.
    is deferred;
    
    MakeVertex (me; V : out TheVertex; P : Pnt from gp)
	---Purpose: Returns in <V> a Vertex built with the point <P>.
    is deferred;
    
    ReverseFace(me; F : in out TheFace)
	---Purpose: Change the orientation of the face.
    is deferred;
    
    AddEdgeVertex(me;
    	    	    E      : in out TheEdge; 
    	    	    V      : in     TheVertex;
		    P      : in     Real;
    	    	    direct : Boolean)
	  ---Purpose: Adds the Vertex <V> in the Edge <E>. <P> is the
	  --          parameter of the vertex on the edge. If <direct>
	  --          is False the Vertex is reversed.
    is deferred;

    AddEdgeVertex(me;
    	    	    E      : in out TheEdge; 
    	    	    V      : in     TheVertex;
		    P1,P2  : in     Real)
	  ---Purpose: Adds the Vertex <V> in the Edge <E>. <P1,P2> are
	  --          the parameters of  the vertex on the  edge.  The
	  --          edge is a closed curve.
    is deferred;

    SetParameters(me;
    	    	    E      : in out TheEdge; 
    	    	    V      : in     TheVertex;
		    P1,P2  : in     Real)
	  ---Purpose: <P1,P2> are the parameters of the  vertex on the
	  --          edge.  The edge is a closed curve.
    is deferred;

    AddWireEdge(me;
    	    	    W      : in out TheWire; 
                    E      : in     TheEdge;
    	    	    direct : Boolean)
	  ---Purpose: Adds the Edge <E> in the  Wire <W>, if direct is
	  --          False the Edge is reversed.
    is deferred;

    AddFaceWire(me;
    	    	    F      : in out TheFace; 
                    W      : in     TheWire)
	  ---Purpose: Adds the Wire <W> in  the Face <F>.
    is deferred;

    AddShellFace(me;
    	    	    Sh     : in out TheShell; 
                    F      : in     TheFace)
	  ---Purpose: Adds the Face <F>  in the Shell <Sh>.
    is deferred;

    CompleteEdge(me; E : in out TheEdge)
	---Purpose: This is called once an edge is completed. It gives
	--          the opportunity to perform any post treatment.
    is deferred;
    
    CompleteWire(me; W : in out TheWire)
	---Purpose: This is called once a wire is  completed. It gives
	--          the opportunity to perform any post treatment.
    is deferred;
    
    CompleteFace(me; F : in out TheFace)
	---Purpose: This is called once a face is  completed. It gives
	--          the opportunity to perform any post treatment.
    is deferred;
    
    CompleteShell(me; S : in out TheShell)
	---Purpose: This is called once a shell is  completed. It gives
	--          the opportunity to perform any post treatment.
    is deferred;
    
end Builder from Primitives;


