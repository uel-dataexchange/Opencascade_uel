-- File:	IGESDimen_ToolWitnessLine.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolWitnessLine  from IGESDimen

    ---Purpose : Tool to work on a WitnessLine. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses WitnessLine from IGESDimen,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolWitnessLine;
    ---Purpose : Returns a ToolWitnessLine, ready to work


    ReadOwnParams (me; ent : mutable WitnessLine;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : WitnessLine;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : WitnessLine;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a WitnessLine <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable WitnessLine) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a WitnessLine
    --           (LineFont forced to Rank = 1, DataType forced to 1)

    DirChecker (me; ent : WitnessLine) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : WitnessLine;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : WitnessLine; entto : mutable WitnessLine;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : WitnessLine;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolWitnessLine;
