-- File:        SurfaceStyleBoundary.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSurfaceStyleBoundary from RWStepVisual

	---Purpose : Read & Write Module for SurfaceStyleBoundary

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SurfaceStyleBoundary from StepVisual,
     EntityIterator from Interface

is

	Create returns RWSurfaceStyleBoundary;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable SurfaceStyleBoundary from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : SurfaceStyleBoundary from StepVisual);

	Share(me; ent : SurfaceStyleBoundary from StepVisual; iter : in out EntityIterator);

end RWSurfaceStyleBoundary;
