-- File:	MDataXtd_GeometryRetrievalDriver.cdl
-- Created:	Wed Nov 19 15:58:25 1997
-- Author:	Denis PASCAL
--		<dp@dingox.paris1.matra-dtv.fr>
-- modified     Sergey Zaritchny
---Copyright:	 Matra Datavision 1997



class GeometryRetrievalDriver from MDataXtd  inherits ARDriver from MDF

	---Purpose: 

uses RRelocationTable from MDF,
     Attribute        from PDF,
     Attribute        from TDF, 
     MessageDriver    from CDM

is


    Create(theMessageDriver : MessageDriver from CDM)  -- Version 0
    returns mutable GeometryRetrievalDriver from MDataXtd;
    

    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type: Geometry from PDataXtd.

    NewEmpty (me)  returns mutable Attribute from TDF;


    Paste(me;
    	  Source     :         Attribute from PDF;
    	  Target     : mutable Attribute from TDF;
    	  RelocTable : RRelocationTable  from MDF);

end GeometryRetrievalDriver;
