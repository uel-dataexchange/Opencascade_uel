-- File:        VectorOrDirection.cdl
-- Created:     Fri Dec  1 11:11:11 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class VectorOrDirection from StepGeom inherits SelectType from StepData

	-- <VectorOrDirection> is an EXPRESS Select Type construct translation.
	-- it gathers : Vector, Direction

uses

	Vector,
	Direction
is

	Create returns VectorOrDirection;
	---Purpose : Returns a VectorOrDirection SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a VectorOrDirection Kind Entity that is :
	--        1 -> Vector
	--        2 -> Direction
	--        0 else

	Vector (me) returns any Vector;
	---Purpose : returns Value as a Vector (Null if another type)

	Direction (me) returns any Direction;
	---Purpose : returns Value as a Direction (Null if another type)


end VectorOrDirection;

