-- File:	StepRepr_NextAssemblyUsageOccurrence.cdl
-- Created:	Mon Jul  3 19:47:51 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class NextAssemblyUsageOccurrence from StepRepr
inherits AssemblyComponentUsage from StepRepr

    ---Purpose: Representation of STEP entity NextAssemblyUsageOccurrence

uses
    HAsciiString from TCollection,
    ProductDefinition from StepBasic

is
    Create returns NextAssemblyUsageOccurrence from StepRepr;
	---Purpose: Empty constructor

end NextAssemblyUsageOccurrence;
