-- File:	Image_GPixelField.cdl
-- Created:	Wed Dec  9 12:22:03 1993
-- Author:	Bertand Lesecq
--		<bbl@sparc3>
---Copyright:	 Matra Datavision 1993

private generic class GPixelField from Image (Item as any)

	---Purpose: The class GPixelField represents bi-dimensionnal arrays 
	--          The range of the index start from 0 .

raises
    RangeError from Standard,
    OutOfRange from Standard,
    OutOfMemory from Standard,
    DimensionMismatch from Standard

is
    
    Create (Width, Height:  Integer from Standard) 
    returns  GPixelField from Image
	---Level: Public
    	---Purpose: Creates an array of lower bound <0><0> and upper
    	--          bound <Width-1><Height-1>.   Range from  Standard  error  is
    	--          raised when <Width-1> is less than <0> or <Height-1> is less
    	--          than <0>.
    raises 
    	RangeError  from Standard,
    	OutOfMemory from Standard;


    Create (Width, Height: Integer from Standard; V : Item) 
    returns  GPixelField from Image
	---Level: Public
    	---Purpose: Creates an array of lower bound <0><0> and upper
    	--          bound <Width-1><Height-1>.   Range from  Standard  error  is
    	--          raised when <Width-1> is less than <0> or <Height-1> is less
    	--          than <0>. The array is initialized with <V>.
    raises
    	RangeError  from Standard,
    	OutOfMemory from Standard;

    Destroy (me : in out )
	---Level: Public
    	---Purpose: Frees   the allocated   area corresponding to  the
    	--          array.   If  the array    was  constructed from  a
    	--          DoubleArray the Destroy doesn't delete the area.
        --          
        ---C++: alias ~
    is static;

    Width (me) returns Integer from Standard
	---Level: Public
    	---Purpose: Return the number of columns of <me>.
    	--          
	---C++: inline
    is static ;

    Height (me) returns Integer from Standard
	---Level: Public
    	---Purpose: Returns the number of rows of <me>.
    	--          
        ---C++: inline
    is static;

    UpperX (me) returns Integer from Standard
	---Level: Public
    	---Purpose:  Returns the upper column number of the array.
    	--          
	---C++: inline
    is static ;

    UpperY (me) returns Integer from Standard
	---Level: Public
    	---Purpose:  Returns the upper row number of the array.
    	--          
	---C++: inline
    is static ;

    SetValue (me : in out; X, Y: Integer from Standard; Value: Item) 
	---Level: Public
    	---Purpose: Sets the element of index <X><Y>
    	--          to <Value>.
	---C++: inline
    raises OutOfRange from Standard
    is static ;

    Value (me; X,Y: Integer from Standard) returns any Item
	---Level: Public
    	---Purpose: Returns the value of the element of index 
        --          <X><Y>
    	--
	---C++: inline
    	---C++: alias operator()
    	---C++: return const &
    raises OutOfRange from Standard
    is static;

    ChangeValue (me: in out; X,Y: Integer from Standard) returns any Item
	---Level: Public
    	---Purpose: Returns the value of the element of index 
        --          <X><Y>
    	--
	---C++: inline
    	---C++: alias operator()
    	---C++: return &
    raises OutOfRange from Standard
    is static;

fields

	myWidth       : Integer from Standard ;
        myHeight      : Integer from Standard ;
	myDeletable   : Boolean;
    	myData        : Address;
	
end GPixelField ;
