-- File:	StepShape_FaceBasedSurfaceModel.cdl
-- Created:	Fri Dec 28 16:02:01 2001 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class FaceBasedSurfaceModel from StepShape
inherits GeometricRepresentationItem from StepGeom

    ---Purpose: Representation of STEP entity FaceBasedSurfaceModel

uses
    HAsciiString from TCollection,
    HArray1OfConnectedFaceSet from StepShape

is
    Create returns FaceBasedSurfaceModel from StepShape;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aFbsmFaces: HArray1OfConnectedFaceSet from StepShape);
	---Purpose: Initialize all fields (own and inherited)

    FbsmFaces (me) returns HArray1OfConnectedFaceSet from StepShape;
	---Purpose: Returns field FbsmFaces
    SetFbsmFaces (me: mutable; FbsmFaces: HArray1OfConnectedFaceSet from StepShape);
	---Purpose: Set field FbsmFaces

fields
    theFbsmFaces: HArray1OfConnectedFaceSet from StepShape;

end FaceBasedSurfaceModel;
