-- File:	RWStepShape_RWPointRepresentation.cdl
-- Created:	Thu Dec 12 15:38:08 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWPointRepresentation from RWStepShape

    ---Purpose: Read & Write tool for PointRepresentation

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    PointRepresentation from StepShape

is
    Create returns RWPointRepresentation from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : PointRepresentation from StepShape);
	---Purpose: Reads PointRepresentation

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: PointRepresentation from StepShape);
	---Purpose: Writes PointRepresentation

    Share (me; ent : PointRepresentation from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWPointRepresentation;
