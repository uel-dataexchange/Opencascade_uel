-- File:        FillAreaStyle.cdl
-- Created:     Mon Dec  4 12:02:27 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWFillAreaStyle from RWStepVisual

	---Purpose : Read & Write Module for FillAreaStyle

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     FillAreaStyle from StepVisual,
     EntityIterator from Interface

is

	Create returns RWFillAreaStyle;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable FillAreaStyle from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : FillAreaStyle from StepVisual);

	Share(me; ent : FillAreaStyle from StepVisual; iter : in out EntityIterator);

end RWFillAreaStyle;
