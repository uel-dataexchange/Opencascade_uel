-- File:        DerivedUnit.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWDerivedUnit from RWStepBasic

	---Purpose : Read & Write Module for DerivedUnit

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     DerivedUnit from StepBasic,
     EntityIterator from Interface

is

	Create returns RWDerivedUnit;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable DerivedUnit from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : DerivedUnit from StepBasic);

	Share(me; ent : DerivedUnit from StepBasic; iter : in out EntityIterator);

end RWDerivedUnit;
