-- File:        BSplineCurveWithKnots.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWBSplineCurveWithKnots from RWStepGeom

	---Purpose : Read & Write Module for BSplineCurveWithKnots
	--           Check added by CKY , 7-OCT-1996

uses Check from Interface, ShareTool from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     BSplineCurveWithKnots from StepGeom,
     EntityIterator from Interface

is

	Create returns RWBSplineCurveWithKnots;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable BSplineCurveWithKnots from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : BSplineCurveWithKnots from StepGeom);

	Share(me; ent : BSplineCurveWithKnots from StepGeom; iter : in out EntityIterator);

    	Check(me; ent : BSplineCurveWithKnots from StepGeom; shares : ShareTool; ach : in out Check);

end RWBSplineCurveWithKnots;
