-- File:	GeomToStep_MakeCurve.cdl
-- Created:	Mon Jun 21 10:14:42 1993
-- Author:	Martine LANGLOIS
--		<mla@mastox>
---Copyright:	 Matra Datavision 1993

class MakeCurve from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          Curve from Geom and the class Curve from StepGeom which
    --          describes a Curve from prostep. As Curve is an 
    --          abstract curve this class an access to the sub-class required.
  
uses Curve from Geom,
     Curve from Geom2d,
     Curve from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( C : Curve from Geom ) returns MakeCurve;

Create ( C : Curve from Geom2d ) returns MakeCurve;

Value (me) returns Curve from StepGeom
    raises NotDone
    is static;
    ---C++: return const&
    
fields

    theCurve : Curve from StepGeom;
    	-- The solution from StepGeom
    	
end MakeCurve;



