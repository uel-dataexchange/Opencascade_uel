-- File:	MakeTranslation.cdl
-- Created:	Mon Sep 28 11:52:25 1992
-- Author:	Remi GILET
--		<reg@sdsun2>
---Copyright:	 Matra Datavision 1992

class MakeTranslation

from GCE2d

    	---Purpose: This class implements elementary construction algorithms for a
    	-- translation in 2D space. The result is a
    	-- Geom2d_Transformation transformation.
    	-- A MakeTranslation object provides a framework for:
    	-- -   defining the construction of the transformation,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the result.

uses Pnt2d          from gp,
     Transformation from Geom2d,
     Vec2d          from gp,
     Real           from Standard
     
is

Create(Vect : Vec2d from gp) returns MakeTranslation;
    	---Purpose: Constructs a translation along the vector Vect.  
    
Create(Point1 : Pnt2d from gp;
       Point2 : Pnt2d from gp) returns MakeTranslation;
    	---Purpose: Constructs a translation along the vector
    	--  (Point1,Point2) defined from the point Point1 to the point Point2.
    
Value(me) returns Transformation from Geom2d
    is static;
       ---C++: return const&
       ---Purpose: Returns the constructed transformation.
    
Operator(me) returns Transformation from Geom2d
    is static;
       ---C++: return const&
       ---C++: alias "Standard_EXPORT operator Handle_Geom2d_Transformation() const;"

fields

    TheTranslation : Transformation from Geom2d;

end MakeTranslation;

