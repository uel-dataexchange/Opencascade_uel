-- File:	BRepClass3d_SClassifier.cdl
-- Created:	Mon Jul 15 17:25:58 1996
-- Author:	Laurent BUCHARD
--		<lbr@cracbox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996



class SClassifier from BRepClass3d
     
     ---Purpose: Provides an algorithm to classify a point in a solid.

uses 
    Pnt     from gp,
    Face    from TopoDS,
    Shape   from TopoDS,
    State   from TopAbs,
    SolidExplorer from BRepClass3d
    
raises
    DomainError from Standard
    
    
    
is 
       
    Create 
    	---Purpose: Empty constructor.
    returns SClassifier from BRepClass3d;
    
    
    Create(S   : in out SolidExplorer from BRepClass3d;
           P   :        Pnt from gp;
	   Tol :        Real from Standard)
    	---Purpose: Constructor to classify the point P with the 
    	--          tolerance Tol on the solid S.
    returns SClassifier from BRepClass3d;
    
    
    Perform(me  : in out;
            S   : in out  SolidExplorer from BRepClass3d;
            P   :         Pnt from gp;
	    Tol :         Real from Standard);
    	---Purpose: Classify the point P with the 
    	--          tolerance Tol on the solid S.
    	--          
    PerformInfinitePoint(me  : in out;
                         S   : in out  SolidExplorer from BRepClass3d;
                         Tol :         Real from Standard);
    	---Purpose: Classify an infinite point with the 
    	--          tolerance Tol on the solid S.

    
    Rejected(me)
    	---Purpose: Returns True if the classification has been 
    	--          computed by rejection. 
    	--          The State is then OUT.
    returns Boolean from Standard;
    
    
    State(me)  returns State  from TopAbs;
    	---Purpose: Returns the result of the classification.
    
    IsOnAFace(me) returns Boolean from Standard;
    	---Purpose: Returns True when the point is a point of a face.
    
    Face(me) 
    	---Purpose: Returns the face used to determine the 
    	--          classification. When the state is ON, this is the 
    	--          face containing the point. 
    	--          
    	--          When Rejected() returns True, Face() has no signification.
    returns Face from TopoDS;

	    
    ForceIn(me: in out) 
    	is protected;
	
    ForceOut(me: in out)
    	is protected;


fields

    myFace         : Face       from TopoDS;
    myState        : Integer    from Standard;  -- 1: Rejected     2: IsOnFace  3: In  4: Out
    
end SClassifier;
