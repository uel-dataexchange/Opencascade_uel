-- File:        AutoDesignGroupedItem.cdl
-- Created:     Fri Dec  1 11:11:10 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class AutoDesignGroupedItem from StepAP214 inherits SelectType from StepData

	-- <AutoDesignGroupedItem> is an EXPRESS Select Type construct translation.
	-- it gathers : AdvancedBrepShapeRepresentation, AnnotationSymbol, CsgRepresentation, FacetedBrepShapeRepresentation, GeometricallyBoundedSurfaceShapeRepresentation, GeometricallyBoundedWireframeShapeRepresentation, ManifoldSurfaceShapeRepresentation, NonManifoldSurfaceShapeRepresentation, RepresentationItem, TemplateInstance
	-- Rev4 adds : CsgShapeRepresentation, Representation, ShapeAspect, ShapeRepresentation
	-- Rev4 removes : AnnotationSymbol, CsgRepresentation, NonManifoldSurfaceShapeRepresentation

uses

	AdvancedBrepShapeRepresentation from StepShape,
	CsgShapeRepresentation from StepShape,
	FacetedBrepShapeRepresentation from StepShape,
	GeometricallyBoundedSurfaceShapeRepresentation from StepShape,
	GeometricallyBoundedWireframeShapeRepresentation from StepShape,
	ManifoldSurfaceShapeRepresentation from StepShape,
	Representation from StepRepr,
	RepresentationItem from StepRepr,
	ShapeAspect from StepRepr,
	ShapeRepresentation from StepShape,
	TemplateInstance from StepVisual
is

	Create returns AutoDesignGroupedItem;
	---Purpose : Returns a AutoDesignGroupedItem SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a AutoDesignGroupedItem Kind Entity that is :
	--        1 -> AdvancedBrepShapeRepresentation
	--        2 -> CsgShapeRepresentation
	--        3 -> FacetedBrepShapeRepresentation
	--        4 -> GeometricallyBoundedSurfaceShapeRepresentation
	--        5 -> GeometricallyBoundedWireframeShapeRepresentation
	--        6 -> ManifoldSurfaceShapeRepresentation
	--        7 -> Representation
	--        8 -> RepresentationItem
	--        9 -> ShapeAspect
	--        10 -> ShapeRepresentation
	--        11 -> TemplateInstance
	--        0 else

	AdvancedBrepShapeRepresentation (me) returns any AdvancedBrepShapeRepresentation;
	---Purpose : returns Value as a AdvancedBrepShapeRepresentation (Null if another type)

	CsgShapeRepresentation (me) returns any CsgShapeRepresentation;
	---Purpose : returns Value as a CsgShapeRepresentation (Null if another type)

	FacetedBrepShapeRepresentation (me) returns any FacetedBrepShapeRepresentation;
	---Purpose : returns Value as a FacetedBrepShapeRepresentation (Null if another type)

	GeometricallyBoundedSurfaceShapeRepresentation (me) returns any GeometricallyBoundedSurfaceShapeRepresentation;
	---Purpose : returns Value as a GeometricallyBoundedSurfaceShapeRepresentation (Null if another type)

	GeometricallyBoundedWireframeShapeRepresentation (me) returns any GeometricallyBoundedWireframeShapeRepresentation;
	---Purpose : returns Value as a GeometricallyBoundedWireframeShapeRepresentation (Null if another type)

	ManifoldSurfaceShapeRepresentation (me) returns any ManifoldSurfaceShapeRepresentation;
	---Purpose : returns Value as a ManifoldSurfaceShapeRepresentation (Null if another type)

	Representation (me) returns any Representation;
	---Purpose : returns Value as a Representation (Null if another type)

	RepresentationItem (me) returns any RepresentationItem;
	---Purpose : returns Value as a RepresentationItem (Null if another type)

	ShapeAspect (me) returns any ShapeAspect;
	---Purpose : returns Value as a ShapeAspect (Null if another type)

	ShapeRepresentation (me) returns any ShapeRepresentation;
	---Purpose : returns Value as a ShapeRepresentation (Null if another type)

	TemplateInstance (me) returns any TemplateInstance;
	---Purpose : returns Value as a TemplateInstance (Null if another type)


end AutoDesignGroupedItem;

