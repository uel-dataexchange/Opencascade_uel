-- File:	RWStepBasic_RWThermodynamicTemperatureUnit.cdl
-- Created:	Thu Dec 12 15:38:09 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWThermodynamicTemperatureUnit from RWStepBasic

    ---Purpose: Read & Write tool for ThermodynamicTemperatureUnit

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ThermodynamicTemperatureUnit from StepBasic

is
    Create returns RWThermodynamicTemperatureUnit from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ThermodynamicTemperatureUnit from StepBasic);
	---Purpose: Reads ThermodynamicTemperatureUnit

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ThermodynamicTemperatureUnit from StepBasic);
	---Purpose: Writes ThermodynamicTemperatureUnit

    Share (me; ent : ThermodynamicTemperatureUnit from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWThermodynamicTemperatureUnit;
