-- File:	RWStepFEA_RWFeaModel3d.cdl
-- Created:	Thu Dec 12 17:51:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFeaModel3d from RWStepFEA

    ---Purpose: Read & Write tool for FeaModel3d

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FeaModel3d from StepFEA

is
    Create returns RWFeaModel3d from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FeaModel3d from StepFEA);
	---Purpose: Reads FeaModel3d

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FeaModel3d from StepFEA);
	---Purpose: Writes FeaModel3d

    Share (me; ent : FeaModel3d from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFeaModel3d;
