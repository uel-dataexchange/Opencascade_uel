-- File:        CartesianTransformationOperator3d.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWCartesianTransformationOperator3d from RWStepGeom

	---Purpose : Read & Write Module for CartesianTransformationOperator3d

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     CartesianTransformationOperator3d from StepGeom,
     EntityIterator from Interface

is

	Create returns RWCartesianTransformationOperator3d;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable CartesianTransformationOperator3d from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : CartesianTransformationOperator3d from StepGeom);

	Share(me; ent : CartesianTransformationOperator3d from StepGeom; iter : in out EntityIterator);

end RWCartesianTransformationOperator3d;
