-- File:	RWStepBasic_RWDocumentRepresentationType.cdl
-- Created:	Wed May 10 15:09:06 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWDocumentRepresentationType from RWStepBasic

    ---Purpose: Read & Write tool for DocumentRepresentationType

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    DocumentRepresentationType from StepBasic

is
    Create returns RWDocumentRepresentationType from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : DocumentRepresentationType from StepBasic);
	---Purpose: Reads DocumentRepresentationType

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: DocumentRepresentationType from StepBasic);
	---Purpose: Writes DocumentRepresentationType

    Share (me; ent : DocumentRepresentationType from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWDocumentRepresentationType;
