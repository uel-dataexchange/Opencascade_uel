-- File:        RepresentationRelationshipWithTransformation.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWRepresentationRelationshipWithTransformation from RWStepRepr

	---Purpose : Read & Write Module for RepresentationRelationshipWithTransformation

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     RepresentationRelationshipWithTransformation from StepRepr,
     EntityIterator from Interface

is

	Create returns RWRepresentationRelationshipWithTransformation;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable RepresentationRelationshipWithTransformation from StepRepr);

	WriteStep (me; SW : in out StepWriter; ent : RepresentationRelationshipWithTransformation from StepRepr);

	Share(me; ent : RepresentationRelationshipWithTransformation from StepRepr; iter : in out EntityIterator);

end RWRepresentationRelationshipWithTransformation;
