-- File:        WeekOfYearAndDayDate.cdl
-- Created:     Mon Dec  4 12:02:33 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWWeekOfYearAndDayDate from RWStepBasic

	---Purpose : Read & Write Module for WeekOfYearAndDayDate

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     WeekOfYearAndDayDate from StepBasic

is

	Create returns RWWeekOfYearAndDayDate;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable WeekOfYearAndDayDate from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : WeekOfYearAndDayDate from StepBasic);

end RWWeekOfYearAndDayDate;
