-- File:	Prs3d_Arrow.cdl
-- Created:	Thu Apr 15 10:20:58 1993
-- Author:	Jean-Louis Frenkel
--		<jlf@phylox>
---Copyright:	 Matra Datavision 1993


class Arrow from Prs3d 
    
inherits Root from Prs3d

	---Purpose: provides class methods to draw an arrow at a given
	--          location, along a given direction and using a given 
	--          angle. 
	
uses
    Pnt from gp,
    Dir from gp,
    PlaneAngle from Quantity,
    Length from Quantity,
    Presentation from Prs3d  

   
is
    Draw(myclass; aPresentation: Presentation from Prs3d;
    	    	  aLocation: Pnt from gp; 
    	    	  aDirection: Dir from gp;
		  anAngle: PlaneAngle from Quantity;
                  aLength: Length from Quantity);
    	---Purpose: Defines the representation of the arrow defined by
    	-- the location point aLocation, the direction
    	-- aDirection and the length aLength.
    	-- The angle anAngle defines the angle of opening of the arrow head.
    	-- The presentation object aPresentation stores the
    	-- information defined in this framework.
        
    Fill(myclass; aPresentation: Presentation from Prs3d;
    	    	  aLocation: Pnt from gp; 
    	    	  aDirection: Dir from gp;
		  anAngle: PlaneAngle from Quantity;
                  aLength: Length from Quantity);
    	---Purpose: Defines the representation of the arrow defined by
    	-- the location point aLocation, the direction vector
    	-- aDirection and the length aLength.
    	-- The angle anAngle defines the angle of opening of
    	-- the arrow head, and the drawer aDrawer specifies
    	-- the display attributes which arrows will have.
    	--  With this syntax, no presentation object is created.
    
end Arrow from Prs3d;
