-- File:	StepShape_ToleranceMethodDefinition.cdl
-- Created:	Tue Apr 24 14:24:28 2001
-- Author:	Christian CAILLET
--		<cky@photox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 2001

class ToleranceMethodDefinition  from StepShape    inherits SelectType  from StepData

    ---Purpose : Added for Dimensional Tolerances

uses
    ToleranceValue from StepShape,
    LimitsAndFits from StepShape

is

    Create returns ToleranceMethodDefinition from StepShape;

    CaseNum (me; ent : Transient) returns Integer;
    ---Purpose : Recognizes a kind of ValueQualifier Select Type :
    --           1 -> ToleranceValue from StepShape
    --           2 -> LimitsAndFits from StepShape

    ToleranceValue (me) returns ToleranceValue from StepShape;
    ---Purpose : Returns Value as ToleranceValue

    LimitsAndFits (me) returns LimitsAndFits from StepShape;
    ---Purpose : Returns Value as LimitsAndFits

end ToleranceMethodDefinition;
