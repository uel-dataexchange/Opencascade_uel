-- File:	RWStepFEA_RWFreedomAndCoefficient.cdl
-- Created:	Sat Dec 14 11:02:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFreedomAndCoefficient from RWStepFEA

    ---Purpose: Read & Write tool for FreedomAndCoefficient

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FreedomAndCoefficient from StepFEA

is
    Create returns RWFreedomAndCoefficient from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FreedomAndCoefficient from StepFEA);
	---Purpose: Reads FreedomAndCoefficient

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FreedomAndCoefficient from StepFEA);
	---Purpose: Writes FreedomAndCoefficient

    Share (me; ent : FreedomAndCoefficient from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFreedomAndCoefficient;
