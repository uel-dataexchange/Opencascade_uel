-- File:	RWStepElement_RWSurfaceSection.cdl
-- Created:	Thu Dec 12 17:29:04 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWSurfaceSection from RWStepElement

    ---Purpose: Read & Write tool for SurfaceSection

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    SurfaceSection from StepElement

is
    Create returns RWSurfaceSection from RWStepElement;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : SurfaceSection from StepElement);
	---Purpose: Reads SurfaceSection

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: SurfaceSection from StepElement);
	---Purpose: Writes SurfaceSection

    Share (me; ent : SurfaceSection from StepElement;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWSurfaceSection;
