-- File:	IGESBasic_ToolGroup.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolGroup  from IGESBasic

    ---Purpose : Tool to work on a Group. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses Group from IGESBasic,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolGroup;
    ---Purpose : Returns a ToolGroup, ready to work


    ReadOwnParams (me; ent : mutable Group;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : Group;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : Group;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a Group <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable Group) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a Group
    --           (Null Elements are removed from list)

    DirChecker (me; ent : Group) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : Group;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : Group; entto : mutable Group;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : Group;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolGroup;
