-- File:	RWStepGeom_RWGeomRepContextAndGlobUnitAssCtxAndGlobUncertaintyAssCtx.cdl
-- Created:	Fri Dec  8 09:28:11 1995
-- Author:	Frederic MAUPAS
--		<fma@anion>
---Copyright:	 Matra Datavision 1995





class RWGeomRepContextAndGlobUnitAssCtxAndGlobUncertaintyAssCtx from RWStepGeom

	---Purpose : Read & Write Module for 
	--           GeomRepContextAndGlobUnitAssCtxAndGlobUncertaintyAssCtx

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     GeomRepContextAndGlobUnitAssCtxAndGlobUncertaintyAssCtx from StepGeom,
     EntityIterator from Interface

is

    Create returns RWGeomRepContextAndGlobUnitAssCtxAndGlobUncertaintyAssCtx;
    
    ReadStep (me; 
   	      data : StepReaderData; 
    	      num : Integer;
              ach : in out Check; 
    	      ent : mutable GeomRepContextAndGlobUnitAssCtxAndGlobUncertaintyAssCtx from StepGeom);

    WriteStep (me; SW : in out StepWriter; 
       	       ent : GeomRepContextAndGlobUnitAssCtxAndGlobUncertaintyAssCtx from StepGeom);

    Share(me; 
    	  ent : GeomRepContextAndGlobUnitAssCtxAndGlobUncertaintyAssCtx from StepGeom; iter : in out EntityIterator);

end RWGeomRepContextAndGlobUnitAssCtxAndGlobUncertaintyAssCtx;
