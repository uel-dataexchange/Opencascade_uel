-- File:	TFace.cdl
-- Created:	Mon Dec 17 11:18:44 1990
-- Author:	Remi Lequette
--		<rle@topsn3>
---Copyright:	 Matra Datavision 1990, 1992



class TFace from PTopoDS inherits TShape from PTopoDS

	---Purpose: A topological  Face.

uses
    ShapeEnum from TopAbs

is
    Create returns mutable TFace from PTopoDS;
	---Purpose: the new TFace covers the whole 2D space.
    ---Level: Internal 
    	
    ShapeType(me) returns ShapeEnum from TopAbs;
    ---Level: Internal 

end TFace;
