-- File:        PresentationRepresentationSelect.cdl
-- Created:     Fri Dec  1 11:11:11 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class PresentationRepresentationSelect from StepVisual inherits SelectType from StepData

	-- <PresentationRepresentationSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : PresentationRepresentation, PresentationSet

uses

	PresentationRepresentation,
	PresentationSet
is

	Create returns PresentationRepresentationSelect;
	---Purpose : Returns a PresentationRepresentationSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a PresentationRepresentationSelect Kind Entity that is :
	--        1 -> PresentationRepresentation
	--        2 -> PresentationSet
	--        0 else

	PresentationRepresentation (me) returns any PresentationRepresentation;
	---Purpose : returns Value as a PresentationRepresentation (Null if another type)

	PresentationSet (me) returns any PresentationSet;
	---Purpose : returns Value as a PresentationSet (Null if another type)


end PresentationRepresentationSelect;

