-- File:	BOP_Area2dBuilder.cdl
-- Created:	Thu Dec 21 17:07:40 1995
-- Author:	Jean Yves LEBEY
--		<jyl@meteox>
---Copyright:	 Matra Datavision 1995

class Area2dBuilder from BOP inherits AreaBuilder from BOP

    ---Purpose:  
    
    -- The algorithm is used to construct Faces from a LoopSet,
    -- where the Loop is the composite topological object of the boundary,
    -- here it is a wire(s) or block(s) of edges.
    -- The LoopSet gives an iteration on Loops.
    -- For each Loop  it indicates if it is on the boundary (wire) or if it
    -- results from  an interference (block of edges).
    -- The result of the algorithm is an iteration on areas.
    -- An area is described by a set of Loops.

uses

    LoopSet        from BOP,
    LoopClassifier from BOP
    
is
    Create returns Area2dBuilder;
    	---Purpose:  
    	--- Empty  Constructor 
    	---
    Create(LS :out LoopSet from BOP;  
    	   LC :out LoopClassifier from BOP;
    	   ForceClass : Boolean from Standard = Standard_False)  
    	returns Area2dBuilder;
    	---Purpose:  
    	--- Creates an  object to build faces on
    	--- the (wires,blocks of edge) of <LS>,  
    	--- using the classifier <LC>.
	---
    InitAreaBuilder(me :out;
    	    	    LS :out LoopSet from BOP;  
    	    	    LC :out LoopClassifier from BOP;
    	    	    ForceClass : Boolean = Standard_False) 
    	is redefined;
    	---Purpose:  
    	--- Initializes the object to find the areas of
    	--- the shapes described by <LS>, 
    	--- using the classifier <LC>.
	---
    
end Area2dBuilder;
