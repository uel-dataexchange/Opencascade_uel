-- File:	StepRepr_SpecifiedHigherUsageOccurrence.cdl
-- Created:	Mon Jul  3 20:13:37 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class SpecifiedHigherUsageOccurrence from StepRepr
inherits AssemblyComponentUsage from StepRepr

    ---Purpose: Representation of STEP entity SpecifiedHigherUsageOccurrence

uses
    HAsciiString from TCollection,
    ProductDefinition from StepBasic,
    AssemblyComponentUsage from StepRepr,
    NextAssemblyUsageOccurrence from StepRepr

is
    Create returns SpecifiedHigherUsageOccurrence from StepRepr;
	---Purpose: Empty constructor

    Init (me: mutable; aProductDefinitionRelationship_Id: HAsciiString from TCollection;
                       aProductDefinitionRelationship_Name: HAsciiString from TCollection;
                       hasProductDefinitionRelationship_Description: Boolean;
                       aProductDefinitionRelationship_Description: HAsciiString from TCollection;
                       aProductDefinitionRelationship_RelatingProductDefinition: ProductDefinition from StepBasic;
                       aProductDefinitionRelationship_RelatedProductDefinition: ProductDefinition from StepBasic;
                       hasAssemblyComponentUsage_ReferenceDesignator: Boolean;
                       aAssemblyComponentUsage_ReferenceDesignator: HAsciiString from TCollection;
                       aUpperUsage: AssemblyComponentUsage from StepRepr;
                       aNextUsage: NextAssemblyUsageOccurrence from StepRepr);
	---Purpose: Initialize all fields (own and inherited)

    UpperUsage (me) returns AssemblyComponentUsage from StepRepr;
	---Purpose: Returns field UpperUsage
    SetUpperUsage (me: mutable; UpperUsage: AssemblyComponentUsage from StepRepr);
	---Purpose: Set field UpperUsage

    NextUsage (me) returns NextAssemblyUsageOccurrence from StepRepr;
	---Purpose: Returns field NextUsage
    SetNextUsage (me: mutable; NextUsage: NextAssemblyUsageOccurrence from StepRepr);
	---Purpose: Set field NextUsage

fields
    theUpperUsage: AssemblyComponentUsage from StepRepr;
    theNextUsage: NextAssemblyUsageOccurrence from StepRepr;

end SpecifiedHigherUsageOccurrence;
