-- File:        RightCircularCylinder.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWRightCircularCylinder from RWStepShape

	---Purpose : Read & Write Module for RightCircularCylinder

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     RightCircularCylinder from StepShape,
     EntityIterator from Interface

is

	Create returns RWRightCircularCylinder;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable RightCircularCylinder from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : RightCircularCylinder from StepShape);

	Share(me; ent : RightCircularCylinder from StepShape; iter : in out EntityIterator);

end RWRightCircularCylinder;
