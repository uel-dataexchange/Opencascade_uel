-- File:	DNaming_CylinderDriver.cdl
-- Created:	Mon May  4 11:31:37 2009
-- Author:	Sergey ZARITCHNY <sergey.zaritchny@opencascade.com> 
---Copyright:	Open CasCade SA 2009


class CylinderDriver from DNaming inherits Driver from TFunction

	---Purpose:  Computes Cylinder function

uses
     Label            from TDF, 
     Logbook          from TFunction,
     Function         from TFunction,
     ExtendedString   from TCollection,
     MakeCylinder     from BRepPrimAPI

is
    Create returns mutable CylinderDriver from DNaming;
    ---Purpose: Constructor

    ---Purpose: validation
    --          ==========

    Validate(me; theLog : in out Logbook from TFunction)
    is redefined;
    ---Purpose: Validates labels of a function in <log>.
    --          In regeneration mode this method must be called (by the
    --          solver) even if the function is not executed, to build
    --          the valid label scope.

    ---Purpose: execution of function
    --          ======================

    MustExecute (me; theLog : Logbook from TFunction)
    ---Purpose: Analyse in <log> if the loaded function must be executed
    --          (i.e.arguments are modified) or not.
    --          If the Function label itself is modified, the function must
    --          be executed.
    returns Boolean from Standard
    is redefined;

    Execute (me; theLog : in out Logbook from TFunction)
    ---Purpose: Execute the function and push in <log> the impacted
    --          labels (see method SetImpacted).
    returns Integer from Standard
    is redefined;
 
    LoadNamingDS(me; theResultLabel : Label from TDF; mkCyl : in out MakeCylinder from BRepPrimAPI)  
    is private; 
     
end CylinderDriver;
