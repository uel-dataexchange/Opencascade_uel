-- File:	IGESSelect_SelectDrawingFrom.cdl
-- Created:	Wed Jun  1 15:53:27 1994
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1994


class SelectDrawingFrom  from IGESSelect  inherits SelectDeduct

    ---Purpose : This selection gets the Drawings attached to its input IGES
    --           entities. They are read through thr Single Views, referenced
    --           in Directory Parts of the entities

uses AsciiString from TCollection, EntityIterator, Graph

raises InterfaceError

is

    Create returns mutable SelectDrawingFrom;
    ---Purpose : Creates a SelectDrawingFrom

    HasUniqueResult (me) returns Boolean  is redefined protected;
    ---Purpose : Returns True, because selection works with a ViewSorter which
    --           gives a unique result

    RootResult (me; G : Graph) returns EntityIterator  raises InterfaceError;
    ---Purpose : Selects the Drawings attached (through Single Views in
    --           Directory Part) to input entities

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns the label, with is "Drawings attached"

end SelectDrawingFrom;

