
-- File:	Graphic2d_Marker.cdl
-- Created:	Jeudi 26 Janvier 1995
-- Author:	CAL
-- Modified: TCL G002A, 28-11-00, new section "inquire methods"
-- SAV 04/07/02 : DrawVertex() redefined.

---Copyright:	Matra Datavision 1995

class Marker from Graphic2d inherits Line from Graphic2d

	---Version:

	---Purpose: The primitive Marker

	---Keywords: Primitive, Marker
	---Warning:
	---References:

uses
	Drawer		from Graphic2d,
	GraphicObject	from Graphic2d,
	Length		from Quantity,
	PlaneAngle	from Quantity, 
	FStream         from Aspect,
	IFStream	from Aspect


raises
	MarkerDefinitionError	from Graphic2d

is
	-------------------------
	-- Category: Constructors
	-------------------------

	Create (aGraphicObject: GraphicObject from Graphic2d;
		X, Y: Length from Quantity)
	returns mutable Marker from Graphic2d;
	---Level: Public
	---Purpose: Creates a pixel point marker at position <X>,<Y>
	---Category: Constructors

	Create (aGraphicObject: GraphicObject from Graphic2d;
		anIndex: Integer from Standard;
		X, Y: Length from Quantity;
		aWidth: Length from Quantity;
		anHeight: Length from Quantity;
		anAngle: PlaneAngle from Quantity = 0.0)
	returns mutable Marker from Graphic2d
	---Level: Public
	---Purpose: Creates the predefined marker index <anIndex> 
	--	    at position <X>,<Y> and size <aWidth>,<aHeight>.
	--	    Angle is measured counterclockwise with 0 radian
	--	    at 3 o'clock.
	---Category: Constructors
	---Trigger: Raises MarkerDefinitionError if the
	--	    marker index is <= 0 or undefined in the MarkMap,
	--          or the marker size <aWidth,anHeight> is null.
	raises MarkerDefinitionError from Graphic2d;

	--------------------------
	-- Category: Draw and Pick
	--------------------------

	Draw (me : mutable; aDrawer: Drawer from Graphic2d)
	is static protected;
	---Level: Internal
	---Purpose: Draws the marker <me>.

	Pick (me : mutable; X, Y: ShortReal from Standard;
		aPrecision: ShortReal from Standard;
		aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard
	is static protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the marker <me> is picked,
	--	    Standard_False if not.
	--  Warning: Checks only if the point <X>, <Y> is in the
	--	    boundary rectangle of <me>

	DrawVertex( me : mutable; aDrawer: Drawer from Graphic2d;
                    anIndex: Integer from Standard)
        is redefined protected;

     --------------------------------------
	-- Category: Inquire methods
	--------------------------------------

    Position( me; X, Y: out Length from Quantity );  
	---Level: Public
	---Purpose: returns the coordinates of the position of the marker
	
    Size( me; aW, aH: out Length from Quantity );  
	---Level: Public
	---Purpose: returns the width and height of the marker
	
	Index( me ) returns Integer from Standard;
	---Level: Public
	---Purpose: returns the index of marker in the map of markers
	
    Angle( me ) returns PlaneAngle from Quantity;
	---Level: Public
	---Purpose: returns the angle of the marker

	----------------------------------------------------------------------

	Save( me; aFStream: in out FStream from Aspect ) is virtual;
--	Retrieve( me; aIFStream: in out IFStream from AIS2D ) is virtual;

fields

	myMarkIndex: Integer from Standard;
	myX:		 ShortReal from Standard;
	myY:		 ShortReal from Standard;
	myWidth:	 ShortReal from Standard;
	myHeight:	 ShortReal from Standard;
	myAngle:	 ShortReal from Standard;

end Marker from Graphic2d;
