-- File:	StepShape_EdgeBasedWireframeShapeRepresentation.cdl
-- Created:	Fri Dec 28 16:02:01 2001 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class EdgeBasedWireframeShapeRepresentation from StepShape
inherits ShapeRepresentation from StepShape

    ---Purpose: Representation of STEP entity EdgeBasedWireframeShapeRepresentation

uses
    HAsciiString from TCollection,
    HArray1OfRepresentationItem from StepRepr,
    RepresentationContext from StepRepr

is
    Create returns EdgeBasedWireframeShapeRepresentation from StepShape;
	---Purpose: Empty constructor

end EdgeBasedWireframeShapeRepresentation;
