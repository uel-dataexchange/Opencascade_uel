-- File:        MechanicalDesignGeometricPresentationArea.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWMechanicalDesignGeometricPresentationArea from RWStepVisual

	---Purpose : Read & Write Module for MechanicalDesignGeometricPresentationArea

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     MechanicalDesignGeometricPresentationArea from StepVisual,
     EntityIterator from Interface

is

	Create returns RWMechanicalDesignGeometricPresentationArea;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable MechanicalDesignGeometricPresentationArea from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : MechanicalDesignGeometricPresentationArea from StepVisual);

	Share(me; ent : MechanicalDesignGeometricPresentationArea from StepVisual; iter : in out EntityIterator);

end RWMechanicalDesignGeometricPresentationArea;
