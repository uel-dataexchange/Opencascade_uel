-- File:	StepBasic_RoleAssociation.cdl
-- Created:	Wed May 10 15:09:08 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RoleAssociation from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity RoleAssociation

uses
    ObjectRole from StepBasic,
    RoleSelect from StepBasic

is
    Create returns RoleAssociation from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aRole: ObjectRole from StepBasic;
                       aItemWithRole: RoleSelect from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Role (me) returns ObjectRole from StepBasic;
	---Purpose: Returns field Role
    SetRole (me: mutable; Role: ObjectRole from StepBasic);
	---Purpose: Set field Role

    ItemWithRole (me) returns RoleSelect from StepBasic;
	---Purpose: Returns field ItemWithRole
    SetItemWithRole (me: mutable; ItemWithRole: RoleSelect from StepBasic);
	---Purpose: Set field ItemWithRole

fields
    theRole: ObjectRole from StepBasic;
    theItemWithRole: RoleSelect from StepBasic;

end RoleAssociation;
