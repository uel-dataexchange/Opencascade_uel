-- File:        TemplateInstance.cdl
-- Created:     Mon Dec  4 12:02:32 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWTemplateInstance from RWStepVisual

	---Purpose : Read & Write Module for TemplateInstance

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     TemplateInstance from StepVisual,
     EntityIterator from Interface

is

	Create returns RWTemplateInstance;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable TemplateInstance from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : TemplateInstance from StepVisual);

	Share(me; ent : TemplateInstance from StepVisual; iter : in out EntityIterator);

end RWTemplateInstance;
