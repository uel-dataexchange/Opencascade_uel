-- File:	StepToGeom_MakeCartesianPoint.cdl
-- Created:	Fri Jun 11 18:43:50 1993
-- Author:	Martine LANGLOIS
---Copyright:	 Matra Datavision 1993

class MakeCartesianPoint from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          CartesianPoint from StepGeom which describes a point from
    --          Prostep and CartesianPoint from Geom.
  
uses 
     CartesianPoint from Geom,
     CartesianPoint from StepGeom
     
is 

    Convert ( myclass; SP : CartesianPoint from StepGeom;
                       CP : out CartesianPoint from Geom )
    returns Boolean from Standard;

end MakeCartesianPoint;
