-- File:        StepShape.cdl
-- Created:     Mon Dec  4 12:02:22 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




package RWStepShape 

uses

	StepData, Interface, TCollection, TColStd, StepShape

is


--class ReadWriteModule;

--class GeneralModule;

class RWAdvancedBrepShapeRepresentation;
class RWAdvancedFace;
class RWBlock;
class RWBooleanResult;
class RWBoxDomain;
class RWBoxedHalfSpace;
class RWBrepWithVoids;
class RWClosedShell;
class RWCompoundShapeRepresentation;
class RWConnectedEdgeSet;
class RWConnectedFaceShapeRepresentation;
class RWConnectedFaceSet;
-- Removed from Rev2 to Rev4 : class RWCsgRepresentation;
class RWCsgShapeRepresentation;
class RWCsgSolid;
class RWDefinitionalRepresentationAndShapeRepresentation; -- abv CAX-IF TRJ4 k1_geo-ac
class RWEdge;
class RWEdgeBasedWireframeModel;
class RWEdgeBasedWireframeShapeRepresentation;
class RWEdgeCurve;
class RWEdgeLoop;
class RWExtrudedAreaSolid;
class RWFace;
class RWFaceBasedSurfaceModel;
class RWFaceBound;
class RWFaceOuterBound;
class RWFaceSurface;
class RWFacetedBrep;
class RWFacetedBrepAndBrepWithVoids; -- Added by FMA
class RWFacetedBrepShapeRepresentation;
class RWGeometricCurveSet;
class RWGeometricSet;
class RWGeometricallyBoundedSurfaceShapeRepresentation;
class RWGeometricallyBoundedWireframeShapeRepresentation;
class RWHalfSpaceSolid;
class RWLoop;
class RWManifoldSolidBrep;
class RWManifoldSurfaceShapeRepresentation;
class RWNonManifoldSurfaceShapeRepresentation;
class RWOpenShell;
class RWOrientedClosedShell;
class RWOrientedEdge;
class RWOrientedFace;
class RWOrientedOpenShell;
class RWOrientedPath;
class RWPath;
class RWPolyLoop;
class RWRevolvedAreaSolid;
class RWRightAngularWedge;
class RWRightCircularCone;
class RWRightCircularCylinder;
class RWShapeRepresentation;
class RWShellBasedSurfaceModel;
class RWSolidModel;
class RWSolidReplica;
class RWSphere;
class RWSweptAreaSolid;
class RWTopologicalRepresentationItem;
class RWTorus;
class RWTransitionalShapeRepresentation;
class RWVertex;
class RWVertexLoop;
class RWVertexPoint;
class RWLoopAndPath;

    --  Added from AP214 CC1 to CC2

class RWContextDependentShapeRepresentation;
class RWShapeDefinitionRepresentation;  -- moved from StepRepr

-- Added from CC2 to DIS
class RWSweptFaceSolid;
class RWExtrudedFaceSolid;
class RWRevolvedFaceSolid;

    -- ABV 18 Apr 00: for dimensions and tolerances (Part 47)
    class RWAngularLocation;
    class RWAngularSize;
    class RWDimensionalCharacteristicRepresentation;
    class RWDimensionalLocation;
    class RWDimensionalLocationWithPath;
    class RWDimensionalSize;
    class RWDimensionalSizeWithPath;
    class RWShapeDimensionRepresentation;

    -- CKY 25 APR 2001 : dim.tol, continued (TR7J)
    class RWLimitsAndFits;
    class RWToleranceValue;
    class RWMeasureQualification;
    class RWPlusMinusTolerance;
    class RWPrecisionQualifier;
    class RWTypeQualifier;

    class RWQualifiedRepresentationItem;
    class RWMeasureRepresentationItemAndQualifiedRepresentationItem;
    
--  Added from AP214 IS to DIS
    
    class RWConnectedFaceSubSet;
    class RWSeamEdge;
    class RWSubedge;
    class RWSubface;
    
--- Added for AP209
    class RWPointRepresentation;

--- added for TR12J (GD&T) 
    class RWShapeRepresentationWithParameters;

	---Package Method ---

--	Init;
	---Purpose: enforced the initialisation of the  libraries

end RWStepShape;
