-- File:        PDataStd_ExtStringList.cdl
-- Created:     May 29 11:40:00 2007
-- Author:      Vlad Romashko
--  	    	<vladislav.romashko@opencascade.com>
-- Copyright:   Open CASCADE

class ExtStringList from PDataStd inherits Attribute from PDF

uses 

    HExtendedString from PCollection,
    HArray1OfExtendedString from PColStd

is

    Create 
    returns mutable ExtStringList from PDataStd;

    Init (me : mutable; 
    	  lower, upper : Integer from Standard);

    SetValue (me: mutable; 
    	      index : Integer from Standard; 
    	      value : HExtendedString from PCollection);

    Value (me;  
    	   index : Integer from Standard) 
    returns HExtendedString from PCollection;

    Lower (me) 
    returns Integer from Standard;      

    Upper (me) 
    returns Integer from Standard;   


fields

    myValue     :  HArray1OfExtendedString from PColStd;


end ExtStringList;
