-- File:	RWStepFEA_RWFeaLinearElasticity.cdl
-- Created:	Thu Dec 12 17:51:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFeaLinearElasticity from RWStepFEA

    ---Purpose: Read & Write tool for FeaLinearElasticity

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FeaLinearElasticity from StepFEA

is
    Create returns RWFeaLinearElasticity from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FeaLinearElasticity from StepFEA);
	---Purpose: Reads FeaLinearElasticity

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FeaLinearElasticity from StepFEA);
	---Purpose: Writes FeaLinearElasticity

    Share (me; ent : FeaLinearElasticity from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFeaLinearElasticity;
