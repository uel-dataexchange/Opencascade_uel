-- File:	RWStepAP214_RWAutoDesignDocumentReference.cdl
-- Created:	Tue Aug  4 13:02:51 1998
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1998


class RWAutoDesignDocumentReference from RWStepAP214

	---Purpose : Read & Write Module for AutoDesignDocumentReference

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     AutoDesignDocumentReference from StepAP214,
     EntityIterator from Interface

is

	Create returns RWAutoDesignDocumentReference;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable AutoDesignDocumentReference from StepAP214);

	WriteStep (me; SW : in out StepWriter; ent : AutoDesignDocumentReference from StepAP214);

	Share(me; ent : AutoDesignDocumentReference from StepAP214; iter : in out EntityIterator);

end RWAutoDesignDocumentReference;
