-- File:        RightCircularCone.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWRightCircularCone from RWStepShape

	---Purpose : Read & Write Module for RightCircularCone

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     RightCircularCone from StepShape,
     EntityIterator from Interface

is

	Create returns RWRightCircularCone;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable RightCircularCone from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : RightCircularCone from StepShape);

	Share(me; ent : RightCircularCone from StepShape; iter : in out EntityIterator);

end RWRightCircularCone;
