-- File:        InvisibilityContext.cdl
-- Created:     Fri Dec  1 11:11:11 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class InvisibilityContext from StepVisual inherits SelectType from StepData

	-- <InvisibilityContext> is an EXPRESS Select Type construct translation.
	-- it gathers : PresentationRepresentation, PresentationSet

uses

	PresentationRepresentation,
	PresentationSet
is

	Create returns InvisibilityContext;
	---Purpose : Returns a InvisibilityContext SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a InvisibilityContext Kind Entity that is :
	--        1 -> PresentationRepresentation
	--        2 -> PresentationSet
	--        0 else

	PresentationRepresentation (me) returns any PresentationRepresentation;
	---Purpose : returns Value as a PresentationRepresentation (Null if another type)

	PresentationSet (me) returns any PresentationSet;
	---Purpose : returns Value as a PresentationSet (Null if another type)


end InvisibilityContext;

