-- File:	StepShape_ConnectedFaceShapeRepresentation.cdl
-- Created:	Fri Dec 28 16:02:00 2001 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class ConnectedFaceShapeRepresentation from StepShape
inherits Representation from StepRepr

    ---Purpose: Representation of STEP entity ConnectedFaceShapeRepresentation

uses
    HAsciiString from TCollection,
    HArray1OfRepresentationItem from StepRepr,
    RepresentationContext from StepRepr

is
    Create returns ConnectedFaceShapeRepresentation from StepShape;
	---Purpose: Empty constructor

end ConnectedFaceShapeRepresentation;
