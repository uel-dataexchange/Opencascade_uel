-- File     : Prs2d_Point.cdl
-- Created  : April  2000
-- Author   : Tanya COOL
---Copyright: Matra Datavision 2000

class Point from Prs2d inherits Line from Graphic2d

  ---Purpose: Constructs presentable and selectable Point. 
  --          It's displayed as a definite type Marker from 
  --          Aspect_TypeOfMarker
  
uses 

  Pnt2d          from gp,
  PlaneAngle     from Quantity,
  Length         from Quantity,
  GraphicObject  from Graphic2d,    
  Drawer         from Graphic2d,
  TypeOfMarker   from Aspect,
  FStream        from Aspect 
    
is
  
  Create( aGO     : GraphicObject from Graphic2d;
          aPnt    : Pnt2d         from gp; 
		  aTOM    : TypeOfMarker  from Aspect;
		  aWSize  : Length        from Quantity = 2.0;
          aHSize  : Length        from Quantity = 2.0;
		  anAngle : PlaneAngle    from Quantity = 0.0  ) 
       returns mutable Point from Prs2d;
  ---Purpose: Initializes the Point defined <aPnt>

  --------------------------
  -- Category: Draw and Pick
  --------------------------

  Draw( me : mutable; aDrawer: Drawer from Graphic2d )
      is static protected;
  ---Level: Internal
  ---Purpose: Draws the angle <me>.

  DrawElement( me : mutable; aDrawer: Drawer from Graphic2d;
                 anIndex: Integer from Standard)
        is redefined protected;
  ---Level: Internal
  ---Purpose: Draws element <anIndex> of the point <me>.

  DrawVertex( me : mutable; aDrawer: Drawer from Graphic2d;
                anIndex: Integer from Standard)
        is redefined protected;
  ---Level: Internal
  ---Purpose: Draws vertex <anIndex> of the point <me>.

  Pick( me: mutable; X, Y      : ShortReal from Standard;
		             aPrecision: ShortReal from Standard;
		             aDrawer   : Drawer from Graphic2d)
	 returns Boolean from Standard is static protected;
  ---Level: Internal
  ---Purpose: Returns Standard_True if the point <me> is picked,
  --	    Standard_False if not.
  
  --------------------------------------------------------------------- 
  ---Category: Modifications of the class properties

  SetPoint( me: mutable; aPnt: Pnt2d from gp );
  ---Level: Public
  ---Purpose: Modifies the Point by redefining location <aPnt>

  SetMarker( me: mutable; aTOM: TypeOfMarker from Aspect );
  ---Level: Public
  ---Purpose: Modifies the Point by redefining type of marker

  SetIndex( me: mutable; anInd: Integer from Standard );
  ---Level: Internal
  ---Purpose: Sets the map index of the marker

  --------------------------------------------------------------------- 
  ---Category: Inquire methods
    
  Point( me ) returns Pnt2d from gp;
  ---Level: Public
  ---Purpose: Returns the location of the Point

  Marker( me ) returns TypeOfMarker from Aspect;
  ---Level: Public
  ---Purpose: Returns the type of marker of the Point

  Save( me; aFStream: in out FStream from Aspect ) is virtual;

fields
	
  myPoint   : Pnt2d        from gp;
  myTOM     : TypeOfMarker from Aspect;
  myIndMark : Integer      from Standard;
  myWSize   : Length       from Quantity;
  myHSize   : Length       from Quantity;
  myAngle   : PlaneAngle   from Quantity;
  
end Point;
