-- File:	RWStepFEA_RWCurveElementInterval.cdl
-- Created:	Thu Dec 12 17:51:04 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWCurveElementInterval from RWStepFEA

    ---Purpose: Read & Write tool for CurveElementInterval

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    CurveElementInterval from StepFEA

is
    Create returns RWCurveElementInterval from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : CurveElementInterval from StepFEA);
	---Purpose: Reads CurveElementInterval

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: CurveElementInterval from StepFEA);
	---Purpose: Writes CurveElementInterval

    Share (me; ent : CurveElementInterval from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWCurveElementInterval;
