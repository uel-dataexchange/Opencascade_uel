-- File:	StepBasic_ProductOrFormationOrDefinition.cdl
-- Created:	Tue Jan 28 12:40:35 2003 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class ProductOrFormationOrDefinition from StepBasic
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type ProductOrFormationOrDefinition

uses
    Product from StepBasic,
    ProductDefinitionFormation from StepBasic,
    ProductDefinition from StepBasic

is
    Create returns ProductOrFormationOrDefinition from StepBasic;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of ProductOrFormationOrDefinition select type
	--          1 -> Product from StepBasic
	--          2 -> ProductDefinitionFormation from StepBasic
	--          3 -> ProductDefinition from StepBasic
	--          0 else

    Product (me) returns Product from StepBasic;
	---Purpose: Returns Value as Product (or Null if another type)

    ProductDefinitionFormation (me) returns ProductDefinitionFormation from StepBasic;
	---Purpose: Returns Value as ProductDefinitionFormation (or Null if another type)

    ProductDefinition (me) returns ProductDefinition from StepBasic;
	---Purpose: Returns Value as ProductDefinition (or Null if another type)

end ProductOrFormationOrDefinition;
