-- File:	RWStepAP214_RWAppliedGroupAssignment.cdl
-- Created:	Wed May 10 15:09:06 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWAppliedGroupAssignment from RWStepAP214

    ---Purpose: Read & Write tool for AppliedGroupAssignment

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    AppliedGroupAssignment from StepAP214

is
    Create returns RWAppliedGroupAssignment from RWStepAP214;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : AppliedGroupAssignment from StepAP214);
	---Purpose: Reads AppliedGroupAssignment

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: AppliedGroupAssignment from StepAP214);
	---Purpose: Writes AppliedGroupAssignment

    Share (me; ent : AppliedGroupAssignment from StepAP214;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWAppliedGroupAssignment;
