-- File:	IGESDimen_ToolLeaderArrow.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolLeaderArrow  from IGESDimen

    ---Purpose : Tool to work on a LeaderArrow. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses LeaderArrow from IGESDimen,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolLeaderArrow;
    ---Purpose : Returns a ToolLeaderArrow, ready to work


    ReadOwnParams (me; ent : mutable LeaderArrow;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : LeaderArrow;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : LeaderArrow;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a LeaderArrow <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : LeaderArrow) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : LeaderArrow;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : LeaderArrow; entto : mutable LeaderArrow;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : LeaderArrow;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolLeaderArrow;
