-- File:	Extrema_GExtPC.cdl
-- Created:	Mon Oct 19 11:55:06 1992
-- Author:	Laurent PAINNOT
--		<lpa@phylox>
---Copyright:	 Matra Datavision 1992

generic class GExtPC from Extrema(
    TheCurve          as any;
    TheCurveTool      as any;
    TheExtPElC        as any;
    ThePoint          as any;
    TheVector         as any;
    ThePOnC           as any;
    TheSequenceOfPOnC as any)
    ---Purpose: It calculates all the distances between  a point and a
    --          curve. The   Algorithm finds the  C2  intervals on the
    --          curve.

uses
    SequenceOfBoolean from TColStd,
    SequenceOfReal    from TColStd,
    CurveType         from GeomAbs
     
raises
    NotDone      from StdFail,
    OutOfRange   from Standard,
    TypeMismatch from Standard


    class EPC    instantiates  GenExtPC      from Extrema
    	(TheCurve,
    	 TheCurveTool,
         ThePOnC,
         ThePoint,
         TheVector);

is
    Create returns GExtPC;
    
    Create(P          : ThePoint;
           C          : TheCurve;
           Uinf, Usup : Real from Standard;
           TolF       : Real from Standard = 1.0e-10)
    	---Purpose: It calculates all the distances.
        --          The function F(u)=distance(P,C(u)) has an extremum
        --          when g(u)=dF/du=0. The algorithm searchs all the
        --          zeros inside the definition range of the curve.
      	--          Zeros are searched between uinf and usup.
      	--          Tol  is used to decide to stop the 
      	--          iterations according to the following condition:
      	--          if n is the number of iterations,
      	--          the algorithm stops when abs(F(Un)-F(Un-1)) < Tol.
    returns GExtPC;

    Create(P    : ThePoint;
           C    : TheCurve;
           TolF : Real from Standard = 1.0e-10)
    	---Purpose: It calculates all the distances.
        --          The function F(u)=distance(P,C(u)) has an extremum
        --          when g(u)=dF/du=0. The algorithm searchs all the
        --          zeros inside the definition range of the curve.
      	--          Tol is used to decide to stop the 
      	--          iterations according to the following condition:
      	--          if n is the number of iterations,
      	--          the algorithm stops when abs(F(Un)-F(Un-1)) < Tol.
    returns GExtPC;
    
    Initialize(me : in out; C          : TheCurve;
                            Uinf, Usup : Real from Standard;
                            TolF       : Real from Standard = 1.0e-10)
    	---Purpose: initializes the fields of the algorithm.
    is static;
    
    Perform(me: in out; P: ThePoint)
    	---Purpose: An exception is raised if the fields have not been
    	--          initialized.
    raises TypeMismatch from Standard
    is static;

    IntervalPerform(me: in out; P: ThePoint)
    is static protected;

    IsDone(me) returns Boolean from Standard
    	---Purpose: True if the distances are found.
    is static;
    
    SquareDistance(me; N: Integer from Standard) returns Real from Standard
    	---Purpose: Returns the value of the <N>th extremum square distance.
    raises NotDone    from StdFail,
    	   OutOfRange from Standard
    is static;
    
    NbExt(me) returns Integer from Standard
    	---Purpose: Returns the number of extremum distances.
    raises NotDone from StdFail
    is static;
    
    IsMin(me; N: Integer from Standard) returns Boolean from Standard
    	---Purpose: Returns True if the <N>th extremum distance is a
    	--          minimum.
    raises NotDone    from StdFail,
    	   OutOfRange from Standard
    is static;
    
    Point(me; N: Integer from Standard) returns ThePOnC
    	---Purpose: Returns the point of the <N>th extremum distance.
    raises NotDone    from StdFail, 
    	   OutOfRange from Standard
    is static;
    
    TrimmedSquareDistances(me; dist1: out Real from Standard;
                         dist2: out Real from Standard;
    	    	    	 P1: out ThePoint;
    	    	    	 P2: out ThePoint)
    	---Purpose: if the curve is a trimmed curve,
    	--          dist1 is a square distance between <P> and the point
    	--          of parameter FirstParameter <P1> and
    	--          dist2 is a square distance between <P> and the point
    	--          of parameter LastParameter <P2>.
    is static;

    
    
fields
    myC:       Address            from Standard;
    Pf:        ThePoint;
    Pl:        ThePoint;
    myExtPElC: TheExtPElC;
    mypoint:   TheSequenceOfPOnC;
    mydone:    Boolean            from Standard;
    mydist1:   Real               from Standard;
    mydist2:   Real               from Standard;
    myExtPC:   EPC                from Extrema;
    mytolu:    Real               from Standard;
    mytolf:    Real               from Standard;
    mysample:  Integer            from Standard;
    myintuinf: Real               from Standard;
    myintusup: Real               from Standard;
    myuinf:    Real               from Standard;
    myusup:    Real               from Standard;
    type:      CurveType          from GeomAbs;
    myismin:   SequenceOfBoolean  from TColStd;
    mySqDist:  SequenceOfReal     from TColStd;
    
end GExtPC;
