-- File:	BOP_Builder.cdl
-- Created:	Thu Mar 29 11:00:59 2001
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2001


deferred  class Builder from BOP 

	---Purpose:  
	
        --  The Root class to perform a Boolean Operations (BO)

uses 

    Shape from TopoDS, 
    Operation from BOP, 
    HistoryCollector from BOP,
    ShapeEnum from TopAbs, 
    DSFiller  from BOPTools,
    PDSFiller from BOPTools, 
     
    IndexedDataMapOfShapeListOfShape from TopTools, 
    ListOfShape       from TopTools, 
    IndexedMapOfShape from TopTools 

--raises

is  

    Initialize 
    	returns Builder from BOP; 
    ---Purpose:  
    --- Empty constructor;
    ---	    
    SetShapes       (me:out; 
    	             aS1: Shape from TopoDS;    	 
    	             aS2: Shape from TopoDS);  
    ---Purpose:  
    --  Set shapes (arguments) to perform BO        
    ---
    SetOperation    (me:out; 
    	    	     anOp:Operation from BOP); 
    ---Purpose:  
    --  Set type of the BO to perform    	     
    -- 
    SetManifoldFlag (me:out; 
                     aFlag:Boolean from Standard);  
    ---Purpose: Set the flag to allow the result  
    --          be manifold or non-manifold (not used) 
    --
    Shape1  (me) 
    	returns Shape from TopoDS; 
    ---C++:  return const &  
    ---Purpose:   
    --  Selector
    --
    Shape2  (me) 
    	returns Shape from TopoDS; 
    ---C++:  return const &   
    ---Purpose:   
    --  Selector
    --
    Operation  (me) 
    	returns Operation from BOP; 
    ---Purpose:   
    --  Selector
    -- 
    ManifoldFlag(me) 
    	returns  Boolean from Standard; 
    ---Purpose:   
    --  Selector
    --	
    IsDone(me) 
    	returns  Boolean  from  Standard ;     	 
    ---Purpose:   
    --	Selector
    -- 
    ErrorStatus (me) 
    	returns  Integer  from  Standard;      	 
    ---Purpose:   
    --  Selector
    --
    Result(me) 
     	returns Shape from TopoDS ;
    ---C++:  return const &  
    ---Purpose:   
    --  Returns the result of the BO      
    -- 
    Do    (me:out) 
    	is virtual;    
    ---Purpose:   
    --           Does the BO from the beggining to the end, 
    --           i.e.  create new DataStructure, DSFiller,         
    --           compute all  interferences, compute states, 
    --           build result etc   
    --
    DoWithFiller  (me:out; 
    	    	   aDSF: DSFiller from BOPTools) 
    	is virtual; 	 
    ---Purpose:   
    --  Does the BO using existing Filler to the end        
    --    
    BuildResult (me:out) 
	is  virtual;	 
    ---Purpose:   
    --  Constructs the final result of the BO 
    --   
    Destroy (me: in out) 
	is  virtual;     
    ---C++: alias "Standard_EXPORT virtual ~BOP_Builder(){Destroy();}" 
    ---Purpose:   
    --  Destructor 
    --     
    SortTypes  (myclass; 
    	    	aType1:out ShapeEnum from TopAbs;  
    	    	aType2:out ShapeEnum from TopAbs);  
    ---Purpose:   
    --  Sort types of shapes as integers in increasing order        
    -- 
    Modified (me;  
    	    	aS : Shape from TopoDS)  
	returns ListOfShape from TopTools; 
    ---C++:  return const & 
    ---Purpose:   
    -- Returns the list  of shapes modified from the shape aS      
    --  
    IsDeleted(me; 
    	    	aS : Shape from TopoDS) 
	returns  Boolean from Standard;  
    ---Purpose:   
    -- Returns TRUE if the result does  not contain the shape aS        
    --   
    FillModified(me:out) 
    	is  protected; 
    ---Purpose:   
    -- Fill the list  of shapes modified from the shape aS.    
    -- For Internal usage 
    --      	     
    FillModified(me:out; 
    	    	aS : Shape from TopoDS; 
    	    	aL : ListOfShape from TopTools) 
	is  protected;	 
    ---Purpose:   
    -- Fill the list  of shapes modified from the shape aS. 
    -- For Internal usage    
    --  
    FillModified(me:out; 
    	    	aE : Shape from TopoDS; 
    	    	aSp: Shape from TopoDS) 
	is  protected;	 
    ---Purpose:   
    -- Fill the list  of shapes modified from the shape aS    
    -- For Internal usage   
    -- 
    SectionEdges (me)  
	returns ListOfShape from TopTools; 
    ---C++:  return const & 
    ---Purpose:   
    -- Returns the list of shapes that are parts of BO "Section" 
    -- for  given arguments. 
    -- For Internal usage       
    --   

    SetHistoryCollector(me: in out; theHistory: HistoryCollector from BOP)
    	is virtual;

    GetHistoryCollector(me)
    	returns HistoryCollector from BOP;

fields 

    myShape1       : Shape from TopoDS      
    	is protected;  
    myShape2       : Shape from TopoDS      
    	is protected;   
    myOperation    : Operation from BOP     
    	is protected; 
    myManifoldFlag : Boolean from Standard  
    	is protected;  	     
    myIsDone       : Boolean from Standard  
    	is protected;      	  
    myErrorStatus  : Integer from Standard  
    	is protected;    
    myResult       : Shape   from TopoDS    
    	is protected;
    myDraw         : Integer   from Standard  
    	is protected; 
    myDSFiller     : PDSFiller from BOPTools  
    	is  protected; 
    myResultMap    : IndexedMapOfShape from TopTools   
    	is  protected; 
    myModifiedMap  : IndexedDataMapOfShapeListOfShape from TopTools   
    	is  protected; 
    myEmptyList    : ListOfShape from TopTools   
    	is  protected;    
    mySectionEdges : ListOfShape from TopTools   
    	is  protected; 

    myHistory: HistoryCollector from BOP
    	is protected;
end Builder;

