-- File:	IGESGraph_ToolTextDisplayTemplate.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolTextDisplayTemplate  from IGESGraph

    ---Purpose : Tool to work on a TextDisplayTemplate. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses TextDisplayTemplate from IGESGraph,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolTextDisplayTemplate;
    ---Purpose : Returns a ToolTextDisplayTemplate, ready to work


    ReadOwnParams (me; ent : mutable TextDisplayTemplate;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : TextDisplayTemplate;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : TextDisplayTemplate;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a TextDisplayTemplate <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : TextDisplayTemplate) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : TextDisplayTemplate;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : TextDisplayTemplate; entto : mutable TextDisplayTemplate;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : TextDisplayTemplate;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolTextDisplayTemplate;
