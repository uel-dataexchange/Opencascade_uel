-- File:	RWStepShape_RWRevolvedFaceSolid.cdl
-- Created:	Mon Mar 15 15:59:48 1999
-- Author:	data exchange team
--		<det@androx.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class RWRevolvedFaceSolid from RWStepShape 

	---Purpose: 

uses
     Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     RevolvedFaceSolid from StepShape,
     EntityIterator from Interface


is
    	Create returns RWRevolvedFaceSolid;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable RevolvedFaceSolid from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : RevolvedFaceSolid from StepShape);

	Share(me; ent : RevolvedFaceSolid from StepShape; iter : in out EntityIterator);



end RWRevolvedFaceSolid;
