-- File:	TopOpeBRep_ShapeIntersector.cdl
-- Created:	Fri May  7 17:03:26 1993
-- Author:	Jean Yves LEBEY
--		<jyl@topsn3>
---Copyright:	 Matra Datavision 1993


class ShapeIntersector from TopOpeBRep

---Purpose: Intersect two shapes.
--          
--          A GeomShape is a  shape with a geometric domain, i.e.
--          a Face or an Edge.
--          
--          The purpose   of  the  ShapeIntersector is   to  find
--          couples  of  intersecting   GeomShape  in  two Shapes
--          (which can   be  any kind of  topologies  : Compound,
--          Solid, Shell, etc... )
--          
--          It  is in charge  of  exploration  of the shapes  and
--          rejection. For this it is provided with two tools :
--            
--            - ShapeExplorer from TopOpeBRepTool.
--            - ShapeScanner from TopOpeBRep which implements bounding boxes.
--
--      Let S1,S2 the shapes sent to InitIntersection(S1,S2) method :
--          - S1 is always SCANNED by a ShapeScanner from TopOpeBRep.
--          - S2 is always EXPLORED by a ShapeExplorer from TopOpeBRepTool.
     
uses

    State from TopAbs,
    Orientation from TopAbs,
    Shape from TopoDS,
    Face from TopoDS,
    HBoxTool from TopOpeBRepTool,
    ShapeTool from TopOpeBRepTool,
    ShapeExplorer from TopOpeBRepTool,
    ShapeScanner from TopOpeBRep,
    FacesIntersector from TopOpeBRep,
    EdgesIntersector from TopOpeBRep,
    FaceEdgeIntersector from TopOpeBRep, 
    --modified by NIZNHY-PKV Fri Sep 24 11:02:16 1999  f
    ListOfShape  from  TopTools 
    --modified by NIZNHY-PKV Fri Sep 24 11:02:19 1999  t
is

    -- -------------------------------
    -- intersection between two shapes
    -- -------------------------------

    Create returns ShapeIntersector from TopOpeBRep;

    InitIntersection(me : in out; S1,S2 : Shape from TopoDS) 
    ---Purpose: Initialize the intersection of shapes S1,S2.
    is static;

    InitIntersection(me : in out; S1,S2 : Shape from TopoDS; 
                                  F1,F2 : Face from TopoDS) 
    ---Purpose: Initialize the intersection of shapes S1,S2.
    is static;

    Reset(me : in out) is static private;
    Init(me : in out; S1,S2 : Shape from TopoDS) is static private;

    Shape(me; Index : Integer from Standard) returns Shape from TopoDS
    ---Purpose: return  the shape  <Index> ( = 1 or 2) given to
    --          InitIntersection().  
    --          Index = 1 will return S1, Index = 2 will return S2.
    ---C++: return const &
    is static;

    MoreIntersection(me) returns Boolean from Standard
    ---Purpose: returns True if there are more intersection
    --          between two the shapes.
    is static;
	
    NextIntersection(me : in out) 
    ---Purpose: search for the next intersection between the two shapes.
    is static;
	
    ChangeFacesIntersector(me : in out) 
    returns FacesIntersector from TopOpeBRep
    ---Purpose: return the current intersection of two Faces.
    ---C++: return &
    is static;

    ChangeEdgesIntersector(me : in out)
    returns EdgesIntersector from TopOpeBRep
    ---Purpose: return the current intersection of two Edges.
    ---C++: return &
    is static;

    ChangeFaceEdgeIntersector(me : in out)
    returns FaceEdgeIntersector from TopOpeBRep
    ---Purpose: return the current intersection of a Face and an Edge.
    ---C++: return &
    is static;

    -- -----------------------------------------
    -- intersection between two geometric shapes
    -- -----------------------------------------
    
    CurrentGeomShape(me; Index : Integer from Standard)  
    returns Shape from TopoDS 
    ---Purpose: return  geometric  shape <Index> ( = 1 or 2 )  of
    --          current intersection.  
    ---C++ : return const &
    is static;

    GetTolerances(me; tol1,tol2 : in out Real from Standard)
    ---Purpose: return  MAX of intersection tolerances with
    --          which FacesIntersector from TopOpeBRep was working.
    is static;


    SetIntersectionDone(me : in out) is static private;

    -- ----------------------------
    -- Faces intersection (private)
    -- ----------------------------
    
    InitFFIntersection(me : in out)
    is static private;
    FindFFIntersection(me : in out)
    is static private;
    MoreFFCouple(me) returns Boolean from Standard 
    is static private;
    NextFFCouple(me : in out) 
    is static private;

    -- ----------------------------
    -- Edges intersection on SameDomain faces (private)
    -- ----------------------------
    
    InitEEFFIntersection(me : in out)
    is static private;
    FindEEFFIntersection(me : in out)
    is static private;
    MoreEEFFCouple(me) returns Boolean from Standard 
    is static private;
    NextEEFFCouple(me : in out) 
    is static private;
	
    -- ----------------------------
    -- Face/Edge intersection (private)
    -- ----------------------------
    
    InitFEIntersection(me : in out)
    is static private;
    FindFEIntersection(me : in out)
    is static private;
    MoreFECouple(me) returns Boolean from Standard 
    is static private;
    NextFECouple(me : in out) 
    is static private;

	
    -- ----------------------------
    -- Edge/Face intersection (private)
    -- ----------------------------
    
    InitEFIntersection(me : in out)
    is static private;
    FindEFIntersection(me : in out)
    is static private;
    MoreEFCouple(me) returns Boolean from Standard 
    is static private;
    NextEFCouple(me : in out) 
    is static private;

    -- ---------------------
    -- Edge/Edge in 2d space (private)
    -- ---------------------

    InitEEIntersection(me : in out)
    is static private;
    FindEEIntersection(me : in out)
    is static private;
    MoreEECouple(me) returns Boolean from Standard 
    is static private;
    NextEECouple(me : in out) 
    is static private;

    -- debug
    DumpCurrent(me; K : Integer from Standard) is static;
    Index(me; K : Integer from Standard) 
    returns Integer from Standard
    is static;
 
--modified by NIZNHY-PKV Fri Sep 24 10:59:59 1999  f 
    RejectedFaces  (me:out;   
                    anObj:Shape  from  TopoDS;   
                    aReference:Shape  from  TopoDS; 
                    aListOfShape:out  ListOfShape  from  TopTools) ;
--modified by NIZNHY-PKV Fri Sep 24 11:00:03 1999  t    

fields

    myShape1 : Shape from TopoDS;
    myShape2 : Shape from TopoDS;
    
    myHBoxTool : HBoxTool from TopOpeBRepTool;
    myFaceExplorer : ShapeExplorer from TopOpeBRepTool;
    myFaceScanner : ShapeScanner from TopOpeBRep;
    myFFIntersector : FacesIntersector from TopOpeBRep;
    myFFSameDomain : Boolean from Standard;
    
    myEdgeExplorer : ShapeExplorer from TopOpeBRepTool;
    myEdgeScanner : ShapeScanner from TopOpeBRep;
    myEEIntersector : EdgesIntersector from TopOpeBRep;
    
    myFEIntersector : FaceEdgeIntersector from TopOpeBRep;

    myEEFace1,myEEFace2 : Face from TopoDS;
    
    myIntersectionDone : Boolean from Standard;
    myTol1 : Real from Standard;
    myTol2 : Real from Standard;

    myFFDone : Boolean from Standard;         
    myEEFFDone : Boolean from Standard;
    myEFDone : Boolean from Standard;
    myFEDone : Boolean from Standard;
    myEEDone : Boolean from Standard;

    myFFInit : Boolean from Standard;         
    myEEFFInit : Boolean from Standard;
    myEFInit : Boolean from Standard;
    myFEInit : Boolean from Standard;
    myEEInit : Boolean from Standard;

end ShapeIntersector from TopOpeBRep;
