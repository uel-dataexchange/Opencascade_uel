-- File:        AutoDesignGroupAssignment.cdl
-- Created:     Fri Dec  1 11:11:14 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class AutoDesignGroupAssignment from StepAP214 

inherits GroupAssignment from StepBasic

uses

	HArray1OfAutoDesignGroupedItem from StepAP214, 
	AutoDesignGroupedItem from StepAP214, 
	Group from StepBasic
is

	Create returns mutable AutoDesignGroupAssignment;
	---Purpose: Returns a AutoDesignGroupAssignment


	Init (me : mutable;
	      aAssignedGroup : mutable Group from StepBasic);

	Init (me : mutable;
	      aAssignedGroup : mutable Group from StepBasic;
	      aItems : mutable HArray1OfAutoDesignGroupedItem from StepAP214) is virtual;

	-- Specific Methods for Field Data Access --

	SetItems(me : mutable; aItems : mutable HArray1OfAutoDesignGroupedItem);
	Items (me) returns mutable HArray1OfAutoDesignGroupedItem;
	ItemsValue (me; num : Integer) returns AutoDesignGroupedItem;
	NbItems (me) returns Integer;

fields

	items : HArray1OfAutoDesignGroupedItem from StepAP214; -- a SelectType

end AutoDesignGroupAssignment;
