-- File:	Circ2dTanOnRad.cdl
-- Created:	Fri Mar 22 11:45:45 1991
-- Author:	Philippe DAUTRY
--		<fid@phobox>
---Copyright:	 Matra Datavision 1991

class Circ2dTanOnRad

from GccAna

	---Purpose: This class implements the algorithms used to 
	--          create a 2d circle tangent to a 2d entity, 
	--          centered on a curv and with a given radius.
	--          The arguments of all construction methods are :
	--             - The qualified element for the tangency constrains 
	--             (QualifiedCirc, QualifiedLin, Points).
	--             - The Center element (circle, line).
	--             - A real Tolerance.
	--          Tolerance is only used in the limits cases.
    	--          For example : 
    	--          We want to create a circle tangent to an OutsideCirc C1
    	--          centered on a line OnLine with a radius Radius and with
    	--          a tolerance Tolerance.
    	--          If we did not use Tolerance it is impossible to 
    	--          find a solution in the the following case : OnLine is 
    	--          outside C1. There is no intersection point between C1
    	--          and OnLine. The distance between the line and the 
    	--          circle is greater than Radius.
    	--          With Tolerance we will give a solution if the 
    	--          distance between C1 and OnLine is lower than or 
    	--          equal Tolerance.

--inherits Storable from Standard

uses Pnt2d           from gp,
     Lin2d           from gp,
     Circ2d          from gp,
     QualifiedCirc   from GccEnt, 
     QualifiedLin    from GccEnt,
     Array1OfReal    from TColStd,
     Array1OfInteger from TColStd,
     Array1OfCirc2d  from TColgp,
     Array1OfPnt2d   from TColgp,
     Position         from GccEnt,
     Array1OfPosition from GccEnt

raises NegativeValue     from Standard,
       OutOfRange        from Standard,
       NotDone           from StdFail,
       BadQualifier      from GccEnt

is

---Category: On a line ................................................

Create(Qualified1 : QualifiedCirc from GccEnt  ;
       OnLine     : Lin2d         from gp      ;
       Radius     : Real          from Standard;
       Tolerance  : Real          from Standard) returns Circ2dTanOnRad 
    ---Purpose: This methods implements the algorithms used to create 
    --          2d Circles tangent to a circle and centered on a 2d Line 
    --          with a given radius.
    --          Tolerance is used to find solution in every limit cases.
    --          For example Tolerance is used in the case of EnclosedCirc when 
    --          Radius-R1+dist is greater Tolerance (dist is the distance 
    --          between the line and the location of the circ, R1 is the 
    --          radius of the circ) because there is no solution.
raises NegativeValue, BadQualifier;
    ---Purpose: raises NegativeValue in case of NegativeRadius.

Create(Qualified1 : QualifiedLin  from GccEnt  ;
       OnLine     : Lin2d         from gp      ;
       Radius     : Real          from Standard;
       Tolerance  : Real          from Standard) returns Circ2dTanOnRad 
    ---Purpose: This methods implements the algorithms used to create 
    --          2d Circles tangent to a 2d Line and centered on a 2d Line 
    --          with a given radius.
    --          Tolerance is used to find solution in every limit cases.
raises NegativeValue, BadQualifier;
    ---Purpose: raises NegativeValue in case of NegativeRadius.

Create(Point1     : Pnt2d         from gp      ;
       OnLine     : Lin2d         from gp      ;
       Radius     : Real          from Standard;
       Tolerance  : Real          from Standard) returns Circ2dTanOnRad 
    ---Purpose: This methods implements the algorithms used to create 
    --          2d Circles passing through a 2d Point and centered on a 
    --          2d Line with a given radius.
    --          Tolerance is used to find solution in every limit cases.
raises NegativeValue;
    -- raises NegativeValue in case of NegativeRadius.

---Category: On a circle ................................................

Create(Qualified1 : QualifiedCirc from GccEnt  ;
       OnCirc     : Circ2d        from gp      ;
       Radius     : Real          from Standard;
       Tolerance  : Real          from Standard) returns Circ2dTanOnRad 
    ---Purpose: This methods implements the algorithms used to create 
    --          2d Circles tangent to a circle and centered on a 2d Circle 
    --          with a given radius.
    --          Tolerance is used to find solution in every limit cases.
raises NegativeValue, BadQualifier;
    ---Purpose: raises NegativeValue in case of NegativeRadius.

Create(Qualified1 : QualifiedLin  from GccEnt  ;
       OnCirc     : Circ2d        from gp      ;
       Radius     : Real          from Standard;
       Tolerance  : Real          from Standard) returns Circ2dTanOnRad 
    ---Purpose: This methods implements the algorithms used to create 
    --          2d Circles tangent to a 2d Line and centered on a 2d Line 
    --          with a given radius.
    --          Tolerance is used to find solution in every limit cases.
raises NegativeValue, BadQualifier;
    ---Purpose: raises NegativeValue in case of NegativeRadius.

Create(Point1     : Pnt2d         from gp      ;
       OnCirc     : Circ2d        from gp      ;
       Radius     : Real          from Standard;
       Tolerance  : Real          from Standard) returns Circ2dTanOnRad 
    ---Purpose: This methods implements the algorithms used to create 
    --          2d Circles passing through a 2d Point and centered on a 
    --          2d Line with a given radius.
    --          Tolerance is used to find solution in every limit cases.
raises NegativeValue;
    ---Purpose: raises NegativeValue in case of NegativeRadius.

-- -- ....................................................................

IsDone(me) returns Boolean from Standard
is static;
    ---Purpose: Returns true if the construction algorithm does not fail
    --          (even if it finds no solution).
    --          Note: IsDone protects against a failure arising from a
    --          more internal intersection algorithm, which has
    --          reached its numeric limits.

NbSolutions(me) returns Integer from Standard
    ---Purpose: This method returns the number of circles, representing solutions.
    --          Raises NotDone if the construction algorithm didn't succeed.
raises NotDone
is static;
    	
ThisSolution(me                           ; 
    	     Index : Integer from Standard) returns Circ2d from gp
    ---Purpose: Returns the solution number Index and raises OutOfRange 
    --   	exception if Index is greater than the number of solutions.
    --          Be careful: the Index is only a way to get all the 
    --          solutions, but is not associated to theses outside the 
    --          context of the algorithm-object.
    -- Raises NotDone if the construction algorithm  didn't succeed.
    --          It raises OutOfRange if Index is greater than the 
    --          number of solutions
raises OutOfRange, NotDone
is static;
       

WhichQualifier(me                                  ;
    	       Index   :     Integer  from Standard;
	       Qualif1 : out Position from GccEnt  )
raises OutOfRange, NotDone
is static;
    ---Purpose: Returns the qualifier Qualif1 of the tangency argument
    --     for the solution of index Index computed by this algorithm.
    --     The returned qualifier is:
    -- -   that specified at the start of construction when the
    --   solutions are defined as enclosed, enclosing or
    --   outside with respect to the argument, or
    -- -   that computed during construction (i.e. enclosed,
    --   enclosing or outside) when the solutions are defined
    --   as unqualified with respect to the argument, or
    -- -   GccEnt_noqualifier if the tangency argument is a point.
    -- Exceptions
    -- Standard_OutOfRange if Index is less than zero or
    -- greater than the number of solutions computed by this algorithm.
    -- StdFail_NotDone if the construction fails. 
        
Tangency1(me                                     ;
          Index         : Integer   from Standard;
          ParSol,ParArg : out Real  from Standard;
          PntSol        : out Pnt2d from gp      )
    ---Purpose: Returns informations about the tangency point between the 
    --          result number Index and the first argument.
    --          ParSol is the intrinsic parameter of the point on the 
    --          solution curv.
    --          ParArg is the intrinsic parameter of the point on the 
    --          argument curv.
    --          PntSol is the tangency point on the solution curv.
    --          PntArg is the tangency point on the argument curv.
    --    Raises NotDone if the construction algorithm didn't succeed.
    --          It raises OutOfRange if Index is greater than the 
    --          number of solutions.
raises OutOfRange, NotDone
is static;
  
CenterOn3 (me                                     ;
           Index         : Integer   from Standard;
           ParArg        : out Real  from Standard;
           PntSol        : out Pnt2d from gp      )
    ---Purpose: Returns informations about the center (on the curv) 
    --          of the result.
    --          ParArg is the intrinsic parameter of the point on 
    --          the argument curv.
    --          PntSol is the center point of the solution curv.
--    Raises NotDone if the construction algorithm  didn't succeed.
    --          It raises OutOfRange if Index is greater than the 
    --          number of solutions.
raises OutOfRange, NotDone
is static;
   

IsTheSame1(me                           ;
           Index : Integer from Standard) returns Boolean from Standard
    ---Purpose: Returns True if the solution number Index is equal to 
    --          the first argument and False in the other cases.
--    Raises NotDone if the construction algorithm  didn't succeed.
    --          It raises OutOfRange if Index is greater than the 
    --          number of solutions.
raises OutOfRange, NotDone
is static;
   

fields

    WellDone : Boolean from Standard;
    ---Purpose: True if the algorithm succeeded.

    NbrSol   : Integer from Standard;
    ---Purpose: The number of possible solutions. We have to decide about the
    --          status of the multiple solutions...

    cirsol   : Array1OfCirc2d from TColgp;
    ---Purpose : The solutions.

    qualifier1 : Array1OfPosition from GccEnt;
    -- The qualifiers of the first argument.

    TheSame1 : Array1OfInteger from TColStd;
    ---Purpose: 1 if the solution and the first argument are the same in the 
    -- tolerance of Tolerance.
    -- 0 in the other cases.

    pnttg1sol   : Array1OfPnt2d from TColgp;
    ---Purpose: The tangency point between the solution and the first 
    --          argument on the solution.

    pntcen3   : Array1OfPnt2d from TColgp;
    ---Purpose: The center point of the solution on the first argument.

    par1sol   : Array1OfReal from TColStd;
    ---Purpose: The parameter of the tangency point between the solution 
    --          and the first argument on thesolution.

    pararg1   : Array1OfReal from TColStd;
    ---Purpose: The parameter of the tangency point between the solution 
    --          and the first argument on the first argument.

    parcen3   : Array1OfReal from TColStd;
    ---Purpose: The parameter of the center point of the solution on the 
    --          second argument.

end Circ2dTanOnRad;

