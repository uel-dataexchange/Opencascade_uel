-- File:	IGESAppli_ToolPWBArtworkStackup.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolPWBArtworkStackup  from IGESAppli

    ---Purpose : Tool to work on a PWBArtworkStackup. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses PWBArtworkStackup from IGESAppli,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolPWBArtworkStackup;
    ---Purpose : Returns a ToolPWBArtworkStackup, ready to work


    ReadOwnParams (me; ent : mutable PWBArtworkStackup;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : PWBArtworkStackup;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : PWBArtworkStackup;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a PWBArtworkStackup <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : PWBArtworkStackup) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : PWBArtworkStackup;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : PWBArtworkStackup; entto : mutable PWBArtworkStackup;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : PWBArtworkStackup;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolPWBArtworkStackup;
