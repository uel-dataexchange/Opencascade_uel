-- File:        AutoDesignNominalDateAssignment.cdl
-- Created:     Fri Dec  1 11:11:14 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class AutoDesignNominalDateAssignment from StepAP214 

inherits DateAssignment from StepBasic 

uses

	HArray1OfAutoDesignDatedItem from StepAP214, 
	AutoDesignDatedItem from StepAP214, 
	Date from StepBasic, 
	DateRole from StepBasic
is

	Create returns mutable AutoDesignNominalDateAssignment;
	---Purpose: Returns a AutoDesignNominalDateAssignment


	Init (me : mutable;
	      aAssignedDate : mutable Date from StepBasic;
	      aRole : mutable DateRole from StepBasic) is redefined;

	Init (me : mutable;
	      aAssignedDate : mutable Date from StepBasic;
	      aRole : mutable DateRole from StepBasic;
	      aItems : mutable HArray1OfAutoDesignDatedItem from StepAP214) is virtual;

	-- Specific Methods for Field Data Access --

	SetItems(me : mutable; aItems : mutable HArray1OfAutoDesignDatedItem);
	Items (me) returns mutable HArray1OfAutoDesignDatedItem;
	ItemsValue (me; num : Integer) returns AutoDesignDatedItem;
	NbItems (me) returns Integer;

fields

	items : HArray1OfAutoDesignDatedItem from StepAP214; -- a SelectType

end AutoDesignNominalDateAssignment;
