-- File:	Geom_Transformation.cdl
-- Created:	Wed Mar 10 10:59:19 1993
-- Author:	JCV
--		<fid@phylox>
-- Copyright:	 Matra Datavision 1993


class Transformation from Geom inherits TShared from MMgt


        ---Purpose : Describes how to construct the following elementary transformations
    	-- - translations,
    	-- - rotations,
    	-- - symmetries,
    	-- - scales.
    	--   The Transformation class can also be used to
    	-- construct complex transformations by combining these
    	-- elementary transformations.
    	-- However, these transformations can never change
    	-- the type of an object. For example, the projection
    	-- transformation can change a circle into an ellipse, and
    	-- therefore change the real type of the object. Such a
    	-- transformation is forbidden in this environment and
    	-- cannot be a Geom_Transformation.
        --  The transformation can be represented as follow :
        --  
        --       V1   V2   V3    T       
        --    | a11  a12  a13   a14 |   | x |      | x'|
        --    | a21  a22  a23   a24 |   | y |      | y'|
        --    | a31  a32  a33   a34 |   | z |   =  | z'|
        --    |  0    0    0     1  |   | 1 |      | 1 |
        --
        --  where {V1, V2, V3} defines the vectorial part of the
        --  transformation and T defines the translation part of 
        --  the transformation.
    	-- Note: Geom_Transformation transformations
    	-- provide the same kind of "geometric" services as
    	-- gp_Trsf ones but have more complex data structures.
    	-- The geometric objects provided by the Geom
    	-- package use gp_Trsf transformations in the syntaxes
    	-- Transform and Transformed.
    	-- Geom_Transformation transformations are used in
    	-- a context where they can be shared by several
    	-- objects contained inside a common data structure.


uses Ax1      from gp, 
     Ax2      from gp, 
     Ax3      from gp, 
     Pnt      from gp, 
     Trsf     from gp,
     TrsfForm from gp,
     Vec      from gp

raises ConstructionError from Standard,
       OutOfRange        from Standard

is


  Create   returns mutable Transformation;
        ---Purpose : Creates an identity transformation.


  Create (T : Trsf)  returns mutable Transformation;
        ---Purpose :  Creates a transient copy of T.


  SetMirror (me : mutable; P : Pnt);
        ---Purpose :
        --  Makes the transformation into a symmetrical transformation
        --  with respect to a point P. 
        --  P is the center of the symmetry.


  SetMirror (me : mutable; A1 : Ax1);
        ---Purpose :
        --  Makes the transformation into a symmetrical transformation
        --  with respect to an axis A1. 
        --  A1 is the center of the axial symmetry.


  SetMirror (me : mutable; A2 : Ax2);
        ---Purpose :
        --  Makes the transformation into a symmetrical transformation
        --  with respect to a plane.  The plane of the symmetry is 
        --  defined with the axis placement A2. It is the plane
        --  (Location, XDirection, YDirection).


  SetRotation (me : mutable; A1 : Ax1; Ang : Real);
        ---Purpose :
        --  Makes the transformation into a rotation.
        --  A1 is the axis rotation and Ang is the angular value
        --  of the rotation in radians.


  SetScale (me : mutable; P : Pnt; S : Real);
        ---Purpose :
        --  Makes the transformation into a scale. P is the center of 
        --  the scale and S is the scaling value.


  SetTransformation (me : mutable; FromSystem1, ToSystem2 : Ax3);
        ---Purpose :
        --  Makes a transformation allowing passage from the coordinate
        --  system "FromSystem1" to the coordinate system "ToSystem2".
        --- Example :
        --  In a C++ implementation :
        --  Real x1, y1, z1;  // are the coordinates of a point in the
        --                    // local system FromSystem1
        --  Real x2, y2, z2;  // are the coordinates of a point in the
        --                    // local system ToSystem2
        --  gp_Pnt P1 (x1, y1, z1) 
        --  Geom_Transformation T;
        --  T.SetTransformation (FromSystem1, ToSystem2);
        --  gp_Pnt P2 = P1.Transformed (T);
        --  P2.Coord (x2, y2, z2);


  SetTransformation (me : mutable; ToSystem : Ax3);
        ---Purpose :
        --  Makes the transformation allowing passage from the basic
        --  coordinate system
        --  {P(0.,0.,0.), VX (1.,0.,0.), VY (0.,1.,0.), VZ (0., 0. ,1.) }
        --  to the local coordinate system defined with the Ax2 ToSystem.
        --  Same utilisation as the previous method. FromSystem1 is
        --  defaulted to the absolute coordinate system.


  SetTranslation (me : mutable; V : Vec);
        ---Purpose :
        --  Makes the transformation into a translation. 
        --  V is the vector of the translation.


  SetTranslation(me : mutable; P1, P2 : Pnt);            
        ---Purpose :
        --  Makes the transformation into a translation from the point
        --  P1 to the point P2.


  SetTrsf (me : mutable; T : Trsf);
        ---Purpose : Converts the gp_Trsf transformation T into this transformation.
      

  IsNegative (me)  returns Boolean;
        ---Purpose : Checks whether this transformation is an indirect
    	-- transformation: returns true if the determinant of the
    	-- matrix of the vectorial part of the transformation is less than 0.
    
  Form (me)  returns TrsfForm;
        ---Purpose : Returns the nature of this transformation as a value
    	-- of the gp_TrsfForm enumeration.
       
                                                      
  ScaleFactor (me)  returns Real;
        ---Purpose :  Returns the scale value of the transformation. 


  Trsf (me)  returns Trsf;
        ---Purpose :
        --  Returns a non transient copy of <me>.
    	---C++: return const&


  Value (me; Row, Col : Integer)   returns Real 
        ---Purpose :
        --  Returns the coefficients of the global matrix of tranformation.
        --  It is a 3 rows X 4 columns matrix.
     raises OutOfRange;
        ---Purpose :
        --  Raised if  Row < 1 or Row > 3  or  Col < 1 or Col > 4



        ---Purpose :
        --  Computes the reverse transformation. 

  Invert (me : mutable)
     raises ConstructionError;
        ---Purpose :
        --  Raised if the the transformation is singular. This means that 
        --  the ScaleFactor is lower or equal to Resolution from 
        --  package gp.


  Inverted (me)    returns mutable Transformation
     raises ConstructionError;
        ---Purpose :
        --  Raised if the the transformation is singular. This means that 
        --  the ScaleFactor is lower or equal to Resolution from 
        --  package gp.





	
  Multiplied (me; Other : Transformation)  returns mutable Transformation;
        ---Purpose :
        --  Computes the transformation composed with Other and <me>.
        --  <me> * Other.
        --  Returns a new transformation


  Multiply (me : mutable; Other : Transformation);
        ---Purpose :
        --  Computes the transformation composed with Other and <me> .
        --  <me> = <me> * Other.


  Power (me : mutable; N : Integer)
        ---Purpose : 
        --  Computes the following composition of transformations
        --  if N > 0  <me> * <me> * .......* <me>.
        --  if N = 0  Identity
        --  if N < 0  <me>.Invert() * .........* <me>.Invert()

     raises ConstructionError;
        ---Purpose :
        --  Raised if N < 0 and if the transformation is not inversible


  Powered (me; N : Integer) returns Transformation
     raises ConstructionError;
        ---Purpose :
        --  Raised if N < 0 and if the transformation is not inversible
 



  PreMultiply (me : mutable; Other : Transformation);
        ---Purpose :
        --  Computes the matrix of the transformation composed with 
        --  <me> and Other.     <me> = Other * <me>


  Transforms (me; X, Y, Z : in out Real);
        ---Purpose :
        --  Applies the transformation <me> to the triplet {X, Y, Z}.



  Copy (me)  returns mutable Transformation;
    	---Purpose: Creates a new object which is a copy of this transformation.    
fields

  gpTrsf : Trsf;

end;
