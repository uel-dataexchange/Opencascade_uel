-- File:	BRepOffsetAPI_MakeThickSolid.cdl
-- Created:	Tue Feb 13 11:00:32 1996
-- Author:	Yves FRICAUD
--		<yfr@stylox>
---Copyright:	 Matra Datavision 1996


class MakeThickSolid from BRepOffsetAPI inherits MakeOffsetShape from BRepOffsetAPI

	---Purpose: Describes functions to build hollowed solids.
    	-- A hollowed solid is built from an initial solid and a set of
    	-- faces on this solid, which are to be removed. The
    	-- remaining faces of the solid become the walls of the
    	-- hollowed solid, their thickness defined at the time of construction.
    	--        the solid is built from an initial
	--          solid  <S> and a  set of  faces {Fi} from  <S>,
	--          builds a   solid  composed  by two shells closed  by
	--          the {Fi}. First shell <SS>   is composed by all
	--          the faces of <S> expected {Fi}.  Second shell is
	--          the offset shell of <SS>.
    	-- A MakeThickSolid object provides a framework for:
    	-- - defining the cross-section of a hollowed solid,
    	-- - implementing the construction algorithm, and
    	-- - consulting the result.
uses

    MakeOffset  from BRepOffset,
    Mode        from BRepOffset,
    Shape       from TopoDS,
    Face        from TopoDS,
    ListOfShape from TopTools,	
    JoinType    from GeomAbs
    
is


    Create returns MakeThickSolid from BRepOffsetAPI;

    
    Create ( S            : Shape       from TopoDS;
    	     ClosingFaces : ListOfShape from TopTools;
             Offset       : Real        from Standard;
	     Tol          : Real        from Standard  ;
	     Mode         : Mode        from BRepOffset = BRepOffset_Skin;
    	     Intersection : Boolean     from Standard   = Standard_False;
	     SelfInter    : Boolean     from Standard   = Standard_False;
             Join         : JoinType    from GeomAbs    = GeomAbs_Arc)
    	---Purpose:  Constructs a hollowed solid from
    	-- the solid S by removing the set of faces ClosingFaces from S, where:
    	--       Offset defines the thickness of the walls. Its sign indicates
    	--   which side of the surface of the solid the hollowed shape is built on;
    	--  - Tol defines the tolerance criterion for coincidence in generated shapes;
    	--  - Mode defines the construction type of parallels applied to free
    	--   edges of shape S. Currently, only one construction type is
    	--   implemented, namely the one where the free edges do not generate
    	--   parallels; this corresponds to the default value BRepOffset_Skin;
    	--   Intersection specifies how the algorithm must work in order to
    	--   limit the parallels to two adjacent shapes:
    	-- - if Intersection is false (default value), the intersection
    	--   is calculated with the parallels to the two adjacent shapes,
    	--  -     if Intersection is true, the intersection is calculated by
    	--   taking account of all parallels generated; this computation
    	--   method is more general as it avoids self-intersections
    	--   generated in the offset shape from features of small dimensions
    	--   on shape S, however this method has not been completely
    	--   implemented and therefore is not recommended for use;
    	--  -     SelfInter tells the algorithm whether a computation to
    	--   eliminate self-intersections needs to be applied to the
    	--   resulting shape. However, as this functionality is not yet
    	--   implemented, you should use the default value (false);
    	--  - Join defines how to fill the holes that may appear between
    	--   parallels to the two adjacent faces. It may take values
    	--   GeomAbs_Arc or GeomAbs_Intersection:
    	-- - if Join is equal to GeomAbs_Arc, then pipes are generated
    	--           between two free edges of two adjacent parallels,
    	--           and spheres are generated on "images" of vertices;
    	--           it is the default value,
    	-- - if Join is equal to GeomAbs_Intersection,
    	--   then the parallels to the two adjacent faces are
    	--   enlarged and intersected, so that there are no free
    	--   edges on parallels to faces.
    	--   Warnings
    	-- Since the algorithm of MakeThickSolid is based on
    	-- MakeOffsetShape algorithm, the warnings are the same as for
    	-- MakeOffsetShape.
    returns MakeThickSolid from BRepOffsetAPI;
    
    Build (me : in out)
    is redefined;
	---Purpose: Builds the resulting shape (redefined from MakeOffsetShape).
	---Level: Public     


    Modified (me: in out; S : Shape from TopoDS)
    	---Purpose: Returns the list  of shapes modified from the shape
    	--          <S>. 
        ---C++: return const & 
        ---Level: Public
    returns ListOfShape from TopTools
    is redefined virtual;


end MakeThickSolid;
