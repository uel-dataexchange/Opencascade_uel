-- File:        MechanicalDesignGeometricPresentationArea.cdl
-- Created:     Fri Dec  1 11:11:22 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class MechanicalDesignGeometricPresentationArea from StepVisual 

inherits PresentationArea from StepVisual 

uses

	HAsciiString from TCollection, 
	HArray1OfRepresentationItem from StepRepr,
	RepresentationContext from StepRepr
is

	Create returns mutable MechanicalDesignGeometricPresentationArea;
	---Purpose: Returns a MechanicalDesignGeometricPresentationArea


end MechanicalDesignGeometricPresentationArea;
