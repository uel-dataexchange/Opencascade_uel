-- File:        BSplineCurve.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWBSplineCurve from RWStepGeom

	---Purpose : Read & Write Module for BSplineCurve

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     BSplineCurve from StepGeom,
     EntityIterator from Interface

is

	Create returns RWBSplineCurve;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable BSplineCurve from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : BSplineCurve from StepGeom);

	Share(me; ent : BSplineCurve from StepGeom; iter : in out EntityIterator);

end RWBSplineCurve;
