-- File:	StepFEA_ElementGroup.cdl
-- Created:	Thu Dec 12 17:51:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class ElementGroup from StepFEA
inherits FeaGroup from StepFEA

    ---Purpose: Representation of STEP entity ElementGroup

uses
    HAsciiString from TCollection,
    FeaModel from StepFEA,
    HArray1OfElementRepresentation from StepFEA

is
    Create returns ElementGroup from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aGroup_Name: HAsciiString from TCollection;
                       aGroup_Description: HAsciiString from TCollection;
                       aFeaGroup_ModelRef: FeaModel from StepFEA;
                       aElements: HArray1OfElementRepresentation from StepFEA);
	---Purpose: Initialize all fields (own and inherited)

    Elements (me) returns HArray1OfElementRepresentation from StepFEA;
	---Purpose: Returns field Elements
    SetElements (me: mutable; Elements: HArray1OfElementRepresentation from StepFEA);
	---Purpose: Set field Elements

fields
    theElements: HArray1OfElementRepresentation from StepFEA;

end ElementGroup;
