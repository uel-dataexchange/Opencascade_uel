-- File:	Lin2dTanPar.cdl
-- Created:	Wed Apr  3 11:10:27 1991
-- Author:	Remi GILET
--		<reg@topsn2>
---Copyright:	 Matra Datavision 1991

class Lin2dTanPar

from GccAna

	---Purpose: This class implements the algorithms used to create 2d 
	--          line tangent to a circle or a point and parallel to 
	--          another line.
        --          The solution has the same orientation as the 
        --          second argument.
    	-- Describes functions for building a 2D line parallel to a line and:
    	-- -   tangential to a circle, or
    	-- -   passing through a point.
    	-- A Lin2dTanPar object provides a framework for:
    	-- -   defining the construction of 2D line(s),
    	-- -   implementing the construction algorithm, and consulting the result(s).

uses   Pnt2d            from gp,
       Lin2d            from gp,
       QualifiedCirc    from GccEnt,
       Array1OfReal     from TColStd,
       Array1OfLin2d    from TColgp,
       Array1OfPnt2d    from TColgp,
       Position         from GccEnt,
       Array1OfPosition from GccEnt

raises OutOfRange        from Standard,
       BadQualifier      from GccEnt,
       NotDone           from StdFail

is

Create (ThePoint   : Pnt2d         from gp;
        Lin1       : Lin2d         from gp) returns Lin2dTanPar;
    	---Purpose: This method implements the algorithms used to create a 2d 
    	--          line passing through a point and parallel to 
    	--          another line.

Create (Qualified1 : QualifiedCirc from GccEnt;
        Lin1       : Lin2d         from gp    ) returns Lin2dTanPar
raises BadQualifier;
    	---Purpose: This method implements the algorithms used to create a 2d 
    	--          line tangent to a circle and parallel to another line.
    	--          It raises BadQualifier in case of EnclosedCirc.
    	-- Exceptions
    	--  GccEnt_BadQualifier if a qualifier is inconsistent with
    	-- the argument it qualifies (for example, enclosed for a circle).


IsDone(me) returns Boolean from Standard
is static;
    	---Purpose : Returns True if the algorithm succeeded.

NbSolutions(me) returns Integer from Standard
    	---Purpose : Returns the number of solutions.
    	-- Raises NotDone if the construction algorithm  didn't succeed.
raises NotDone
is static;

ThisSolution(me                                  ;
             Index        : Integer from Standard) returns Lin2d 
    	---Purpose : Returns the solution number Index and raises OutOfRange 
    	--           exception if Index is greater than the number of solutions.
    	--           Be careful: the Index is only a way to get all the 
    	--           solutions, but is not associated to those outside the 
    	--           context of the algorithm-object.
    	-- raises NotDone if the construction algorithm 
    	--          didn't succeed.
    	--          It raises OutOfRange if Index is greater than the 
    	--          number of solutions.

raises OutOfRange, NotDone
is static;
   
WhichQualifier(me                                  ;
    	       Index   :     Integer  from Standard;
	       Qualif1 : out Position from GccEnt  )
raises OutOfRange, NotDone
is static;
    	---Purpose: Returns the informations about the qualifiers of the 
    	--          tangency arguments concerning the solution number Index.
    	--          It returns the real qualifiers (the qualifiers given to the 
    	--          constructor method in case of enclosed, enclosing and outside 
    	--          and the qualifiers computed in case of unqualified).
    	-- Raises NotDone if the construction algorithm 
    	--          didn't succeed.
    	--          It raises OutOfRange if Index is greater than the 
    	--          number of solutions.

Tangency1(me                                      ; 
          Index         : Integer    from Standard; 
          ParSol,ParArg : out Real   from Standard;
          Pnt           : out Pnt2d  from gp      )
    	---Purpose : Returns informations about the tangency point between the 
    	--           result number Index and the first argument.
    	--           ParSol is the intrinsic parameter of the point on the 
    	--           solution curv.
    	--           ParArg is the intrinsic parameter of the point on the
    	--           argument curv.
    	--           ParArg is equal 0 when the solution is passing thrue 
    	--           a point. Raises NotDone if the construction algorithm 
    	--          didn't succeed.
    	--          It raises OutOfRange if Index is greater than the 
    	--          number of solutions.
raises OutOfRange, NotDone
is static;
   
fields

    WellDone : Boolean from Standard;
    	---Purpose: True if the algorithm succeeded.

    NbrSol   : Integer from Standard;
    	---Purpose : The number of possible solutions. We have to decide 
    	--           about the status of the multiple solutions...

    linsol   : Array1OfLin2d from TColgp;
    	---Purpose: The solutions.

    qualifier1 : Array1OfPosition from GccEnt;
    	---Purpose: The qualifiers of the first argument.

    pnttg1sol   : Array1OfPnt2d from TColgp;
    	---Purpose: The tangency point between the solution and the 
    	--          first argument on the solution.

    par1sol   : Array1OfReal from TColStd;
    	---Purpose: The parameter of the tangency point between the 
    	--          solution and the first argument on the solution.

    pararg1   : Array1OfReal from TColStd;
    	---Purpose: The parameter of the tangency point between the 
    	--          solution and the first argument on the first argument.

end Lin2dTanPar;

