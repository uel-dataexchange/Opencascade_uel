-- File:	RWStepShape_RWDimensionalCharacteristicRepresentation.cdl
-- Created:	Tue Apr 18 16:42:58 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWDimensionalCharacteristicRepresentation from RWStepShape

    ---Purpose: Read & Write tool for DimensionalCharacteristicRepresentation

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    DimensionalCharacteristicRepresentation from StepShape

is
    Create returns RWDimensionalCharacteristicRepresentation from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : DimensionalCharacteristicRepresentation from StepShape);
	---Purpose: Reads DimensionalCharacteristicRepresentation

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: DimensionalCharacteristicRepresentation from StepShape);
	---Purpose: Writes DimensionalCharacteristicRepresentation

    Share (me; ent : DimensionalCharacteristicRepresentation from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWDimensionalCharacteristicRepresentation;
