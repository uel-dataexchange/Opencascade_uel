-- File:	Vrml_Coordinate3.cdl
-- Created:	Wed Feb  5 13:25:06 1997
-- Author:	Alexander BRIVIN and Dmitry TARASOV
--		<brivin@minox.nizhny.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


class Coordinate3 from Vrml inherits  TShared  from  MMgt

	---Purpose: defines a Coordinate3 node of VRML specifying
	--          properties of geometry and its appearance. 
    	--  This node defines a set of 3D coordinates to be used by a subsequent IndexedFaceSet,  
    	--  IndexedLineSet, or PointSet node. This node does not produce a visible result  
    	--  during rendering; it simply replaces the current coordinates in the rendering  
    	--  state for subsequent nodes to use. 
uses
 
     HArray1OfVec  from  TColgp 

is
    Create ( aPoint : HArray1OfVec  from  TColgp )
    	returns mutable Coordinate3 from Vrml; 
     
    Create  returns mutable Coordinate3 from Vrml;
    
    SetPoint ( me  :  mutable; aPoint : HArray1OfVec  from  TColgp );
    Point ( me )  returns  HArray1OfVec  from  TColgp; 
    
    Print  ( me;  anOStream: in out OStream from Standard) returns OStream from Standard;
    ---C++:  return  & 

fields

    myPoint  : HArray1OfVec  from  TColgp;  -- Coordinate point(s)

end Coordinate3;
