-- File:	StepAP203_CcDesignCertification.cdl
-- Created:	Fri Nov 26 16:26:31 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class CcDesignCertification from StepAP203
inherits CertificationAssignment from StepBasic

    ---Purpose: Representation of STEP entity CcDesignCertification

uses
    Certification from StepBasic,
    HArray1OfCertifiedItem from StepAP203

is
    Create returns CcDesignCertification from StepAP203;
	---Purpose: Empty constructor

    Init (me: mutable; aCertificationAssignment_AssignedCertification: Certification from StepBasic;
                       aItems: HArray1OfCertifiedItem from StepAP203);
	---Purpose: Initialize all fields (own and inherited)

    Items (me) returns HArray1OfCertifiedItem from StepAP203;
	---Purpose: Returns field Items
    SetItems (me: mutable; Items: HArray1OfCertifiedItem from StepAP203);
	---Purpose: Set field Items

fields
    theItems: HArray1OfCertifiedItem from StepAP203;

end CcDesignCertification;
