-- File:        AlienImage_BMPAlienImage.cdl
-- Created:     20/10/98
-- Author:      DCB
---Copyright:   Matravision 1993

class BMPAlienImage from AlienImage inherits AlienUserImage from AlienImage

uses
  BMPAlienData            from AlienImage,
  File                    from OSD,
  AsciiString             from TCollection,
  Image                   from Image

is
  Create
  returns mutable BMPAlienImage from AlienImage;

  Clear( me : in out mutable) ;
  ---Level: Public
  ---Purpose: Frees memory allocated by BMPAlienImage
  ---C++: alias ~

  SetName( me : in out mutable;
           aName : in AsciiString from TCollection) ;
  ---Level: Public
  ---Purpose: Set Image name .

  Name( me : in immutable ) returns AsciiString from TCollection ;
  ---C++: return const &
  ---Level: Public
  ---Purpose: get Image name .

  ToImage( me : in immutable ) 
  returns mutable Image from Image ;
  ---Level: Public
  ---Purpose : convert a BMPAlienImage object to a Image object.

  FromImage( me : in out mutable ; anImage : in Image from Image ) ;
  ---Level: Public
  ---Purpose : convert a Image object to a BMPAlienImage object.

  Read ( me : in out mutable; afile : in out File from OSD )
    returns Boolean from Standard ;
  ---Level: Public
  ---Purpose: Read content of a  BMPAlienImage object from a file .
  --          Returns True if file is a BMP file .

  Write( me : in immutable; afile : in out File from OSD )
  returns Boolean from Standard ;
  ---Level: Public
  ---Purpose: Write content of a  BMPAlienImage object to a file .

fields
  myData : BMPAlienData from AlienImage;

end;
 
