-- File:	STEPConstruct_AP203Context.cdl
-- Created:	Thu Nov 18 19:46:52 1999
-- Author:	Andrey BETENEV
--		<abv@doomox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class AP203Context from STEPConstruct 

    ---Purpose: Maintains context specific for AP203 (required data and
    --          management information such as persons, dates, approvals etc.)
    --          It contains static entities (which can be shared), default
    --          values for person and organisation, and also provides
    --          tool for creating management entities around specific part (SDR).

uses
    Approval from StepBasic,
    DateAndTime from StepBasic,
    PersonAndOrganization from StepBasic,
    SecurityClassificationLevel from StepBasic,
    PersonAndOrganizationRole from StepBasic,
    DateTimeRole from StepBasic,
    ApprovalRole from StepBasic,
    CcDesignPersonAndOrganizationAssignment from StepAP203,
    CcDesignSecurityClassification from StepAP203,
    CcDesignDateAndTimeAssignment from StepAP203,
    CcDesignApproval from StepAP203,
    ApprovalPersonOrganization from StepBasic,
    ApprovalDateTime from StepBasic,
    ShapeDefinitionRepresentation from StepShape,
    NextAssemblyUsageOccurrence from StepRepr,
    ProductCategoryRelationship from StepBasic,
    Part from STEPConstruct

is
    Create returns AP203Context from STEPConstruct;
    	---Purpose: Creates tool and fills constant fields
	    
    --- Entities shared by others by default
	    
    DefaultApproval (me: in out) returns Approval from StepBasic;
    	---Purpose: Returns default approval entity which 
        --          is used when no other data are available    
    SetDefaultApproval (me: in out; app: Approval from StepBasic);
    	---Purpose: Sets default approval
    
    DefaultDateAndTime (me: in out) returns DateAndTime from StepBasic;
    	---Purpose: Returns default date_and_time entity which 
        --          is used when no other data are available
    SetDefaultDateAndTime (me: in out; dt: DateAndTime from StepBasic);
    	---Purpose: Sets default date_and_time entity 
    
    DefaultPersonAndOrganization (me: in out) returns PersonAndOrganization from StepBasic;
    	---Purpose: Returns default person_and_organization entity which 
        --          is used when no other data are available
    SetDefaultPersonAndOrganization (me: in out; po: PersonAndOrganization from StepBasic);
    	---Purpose: Sets default person_and_organization entity 
    
    DefaultSecurityClassificationLevel (me: in out) returns SecurityClassificationLevel from StepBasic;
    	---Purpose: Returns default security_classification_level entity which 
        --          is used when no other data are available
    SetDefaultSecurityClassificationLevel (me: in out; sc: SecurityClassificationLevel from StepBasic);
    	---Purpose: Sets default security_classification_level
    
    RoleCreator (me) returns PersonAndOrganizationRole from StepBasic;
    RoleDesignOwner (me) returns PersonAndOrganizationRole from StepBasic;
    RoleDesignSupplier (me) returns PersonAndOrganizationRole from StepBasic;
    RoleClassificationOfficer (me) returns PersonAndOrganizationRole from StepBasic;
    RoleCreationDate (me) returns DateTimeRole from StepBasic;
    RoleClassificationDate (me) returns DateTimeRole from StepBasic;
    RoleApprover (me) returns ApprovalRole from StepBasic;
    	---Purpose: Return predefined PersonAndOrganizationRole and DateTimeRole 
	--          entities named 'creator', 'design owner', 'design supplier',
	--          'classification officer', 'creation date', 'classification date',
	--          'approver'

    --- Entities instantiated for each part
    
    Init (me: in out; sdr: ShapeDefinitionRepresentation from StepShape);
    	---Purpose: Takes SDR (part) which brings all standard data around part 
	--          (common for AP203 and AP214) and creates all the additional 
	--          entities required for AP203
    
    Init (me: in out; SDRTool: Part from STEPConstruct);
    	---Purpose: Takes tool which describes standard data around part 
	--          (common for AP203 and AP214) and creates all the additional 
	--          entities required for AP203
	--
	--          The created entities can be obtained by calls to methods
        --          GetCreator(), GetDesignOwner(), GetDesignSupplier(), 
        --          GetClassificationOfficer(), GetSecurity(), GetCreationDate(), 
        --          GetClassificationDate(), GetApproval(), 
        --          GetApprover(), GetApprovalDateTime(),
	--          GetProductCategoryRelationship()
    
    Init (me: in out; nauo: NextAssemblyUsageOccurrence from StepRepr);
    	---Purpose: Takes NAUO which describes assembly link to component
	--          and creates the security_classification entity associated to 
        --          it as required by the AP203
	--          
	--          Instantiated (or existing previously) entities concerned
	--          can be obtained by calls to methods
        --          GetClassificationOfficer(), GetSecurity(), 
        --          GetClassificationDate(), GetApproval(), 
        --          GetApprover(), GetApprovalDateTime()
    
--    Init (me: in out; SDRTool: Part from STEPConstruct; 
--                      Model: InterfaceModel from Interface);
    	---Purpose: Takes tool which describes standard data around part 
	--          (common for AP203 and AP214) and takes from model (or creates
        --          if missing) all the additional entities required by AP203

    GetCreator (me) returns CcDesignPersonAndOrganizationAssignment from StepAP203;
    GetDesignOwner (me) returns CcDesignPersonAndOrganizationAssignment from StepAP203;
    GetDesignSupplier (me) returns CcDesignPersonAndOrganizationAssignment from StepAP203;
    GetClassificationOfficer (me) returns CcDesignPersonAndOrganizationAssignment from StepAP203;
    GetSecurity (me) returns CcDesignSecurityClassification from StepAP203;
    GetCreationDate (me) returns CcDesignDateAndTimeAssignment from StepAP203;
    GetClassificationDate (me) returns CcDesignDateAndTimeAssignment from StepAP203;
    GetApproval (me) returns CcDesignApproval from StepAP203;
    GetApprover (me) returns ApprovalPersonOrganization from StepBasic;
    GetApprovalDateTime (me) returns ApprovalDateTime from StepBasic;
    GetProductCategoryRelationship (me) returns ProductCategoryRelationship from StepBasic;
    	---Purpose: Return entities (roots) instantiated for the part by method Init
    
    --- Advanced (rather internal) methods
    
    Clear (me: in out);
    	---Purpose: Clears all fields describing entities specific to each part
	
    InitRoles (me: in out);
    	---Purpose: Initializes constant fields (shared entities)

    InitPart (me: in out; SDRTool: Part from STEPConstruct) is private;
    	---Purpose: Initializes all missing data which are required for part

    InitAssembly (me: in out; nauo: NextAssemblyUsageOccurrence from StepRepr);
    	---Purpose: Initializes all missing data which are required for assembly
	
    InitSecurityRequisites (me: in out);
    	---Purpose: Initializes ClassificationOfficer and ClassificationDate
	--          entities according to Security entity

    InitApprovalRequisites (me: in out);
    	---Purpose: Initializes Approver and ApprovalDateTime
	--          entities according to Approval entity
    
fields

    -- default values (to be replaced by some meaningful externally)
    defApproval              : Approval from StepBasic;
    defDateAndTime           : DateAndTime from StepBasic;
    defPersonAndOrganization : PersonAndOrganization from StepBasic;
    defSecurityClassificationLevel: SecurityClassificationLevel from StepBasic;
    
    -- predefined roles
    roleCreator              : PersonAndOrganizationRole from StepBasic;
    roleDesignOwner          : PersonAndOrganizationRole from StepBasic;
    roleDesignSupplier       : PersonAndOrganizationRole from StepBasic;
    roleClassificationOfficer: PersonAndOrganizationRole from StepBasic;
    roleCreationDate         : DateTimeRole from StepBasic;
    roleClassificationDate   : DateTimeRole from StepBasic;
    roleApprover             : ApprovalRole from StepBasic;

    -- entities created for each part (roots)
    myCreator                : CcDesignPersonAndOrganizationAssignment from StepAP203;
    myDesignOwner            : CcDesignPersonAndOrganizationAssignment from StepAP203;
    myDesignSupplier         : CcDesignPersonAndOrganizationAssignment from StepAP203;
    myClassificationOfficer  : CcDesignPersonAndOrganizationAssignment from StepAP203;
    mySecurity               : CcDesignSecurityClassification from StepAP203;
    myCreationDate           : CcDesignDateAndTimeAssignment from StepAP203;
    myClassificationDate     : CcDesignDateAndTimeAssignment from StepAP203;
    myApproval               : CcDesignApproval from StepAP203;

    myApprover               : ApprovalPersonOrganization from StepBasic;
    myApprovalDateTime       : ApprovalDateTime from StepBasic;
    
    myProductCategoryRelationship: ProductCategoryRelationship from StepBasic;

end AP203Context;
