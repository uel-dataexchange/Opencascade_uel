-- File:	StepToGeom_MakeEllipse2d.cdl
-- Created:	Thu Sep  1 13:56:44 1994
-- Author:	Frederic MAUPAS
---Copyright:	 Matra Datavision 1994

class MakeEllipse2d from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          Ellipse from StepGeom which describes a Ellipse from
    --          Prostep and Ellipse from Geom2d.
  
uses 
     Ellipse from Geom2d,
     Ellipse from StepGeom
     
is 

    Convert ( myclass; SC : Ellipse from StepGeom;
                       CC : out Ellipse from Geom2d )
    returns Boolean from Standard;

end MakeEllipse2d;
