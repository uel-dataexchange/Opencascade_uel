-- File:	GeomFill_BSplineCurves.cdl
-- Created:	Wed Oct  6 10:50:12 1993
-- Author:	Bruno DUMORTIER
--		<dub@sdsun1>
---Copyright:	 Matra Datavision 1993

class BSplineCurves from GeomFill

	---Purpose: An algorithm for constructing a BSpline surface filled
    	-- from contiguous BSpline curves which form its boundaries.
    	-- The algorithm accepts two, three or four BSpline
    	-- curves as the boundaries of the target surface.
    	-- A range of filling styles - more or less rounded, more
    	-- or less flat - is available.
    	-- A BSplineCurves object provides a framework for:
    	-- -   defining the boundaries, and the filling style of the surface
    	-- -   implementing the construction algorithm
    	-- -   consulting the result.
    	-- Warning
    	-- Some problems may show up with rational curves.

uses
    BSplineCurve    from Geom,
    BSplineSurface  from Geom,
    FillingStyle   from GeomFill

raises
    ConstructionError from Standard
is
    Create;
    	---Purpose: Constructs a default BSpline surface framework.
    
    Create( C1, C2, C3, C4 : BSplineCurve  from Geom;
    	    Type           : FillingStyle from GeomFill)
    returns BSplineCurves from GeomFill;
    
    Create( C1, C2, C3 : BSplineCurve  from Geom;
    	    Type       : FillingStyle from GeomFill)
    returns BSplineCurves from GeomFill;
    
    Create( C1, C2 : BSplineCurve  from Geom;
    	    Type   : FillingStyle from GeomFill)
    returns BSplineCurves from GeomFill;
    	---Purpose: Constructs a framework for building a BSpline surface from either
    	-- -   the four contiguous BSpline curves, C1, C2, C3 and C4, or
    	-- -   the three contiguous BSpline curves, C1, C2 and C3, or
    	-- -   the two contiguous BSpline curves, C1 and C2.
    	-- The type of filling style Type to be used is one of:
    	-- -   GeomFill_Stretch - the style with the flattest patch
    	-- -   GeomFill_Coons - a rounded style of patch with
    	--   less depth than that of Curved
    	-- -   GeomFill_Curved - the style with the most rounded
    	--   patch.Constructs a framework for building a BSpline
    	--   surface common to the two BSpline curves, C1 and C2.
    	-- Exceptions
    	-- Standard_ConstructionError if the curves are not contiguous.
    
    Init( me : in out;
    	  C1, C2, C3, C4 : BSplineCurve  from Geom;
    	  Type           : FillingStyle from GeomFill)
    raises
    	ConstructionError from Standard
	---Purpose: if the curves cannot be joined
    is static;
    
    Init( me : in out;
          C1, C2, C3 : BSplineCurve  from  Geom;
    	  Type       : FillingStyle from GeomFill)
    raises
    	ConstructionError from Standard
	---Purpose: if the curves cannot be joined
    is static;
    
    Init( me : in out;
          C1, C2 : BSplineCurve  from  Geom;
    	  Type   : FillingStyle from GeomFill)
    is static;
    	---Purpose: Initializes or reinitializes this algorithm with two, three,
    	-- or four curves - C1, C2, C3, and C4 - and Type, one
    	-- of the following filling styles:
    	-- -   GeomFill_Stretch - the style with the flattest patch
    	-- -   GeomFill_Coons - a rounded style of patch with
    	--   less depth than that of Curved
    	-- -   GeomFill_Curved - the style with the most rounded patch.
    	--   Exceptions
    	-- Standard_ConstructionError if the curves are not contiguous.
        
    Surface(me) returns BSplineSurface from Geom
    	---Purpose: Returns the BSpline surface Surface resulting from
    	-- the computation performed by this algorithm.
    	---C++: return const&
    	---C++: inline
        
    is static;
    
fields

    mySurface : BSplineSurface from Geom;
    
end BSplineCurves;
