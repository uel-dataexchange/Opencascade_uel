-- File:	LocOpe_RevolutionForm.cdl
-- Created:	Mon Oct 20 09:11:01 1997
-- Author:	Olga KOULECHOVA
--		<opt@cleox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997

class RevolutionForm from LocOpe 

	---Purpose: Defines a revolution form (using Revol from BRepSweep)
	--     with modifications provided for the RevolutionForm feature.
uses DataMapOfShapeListOfShape from TopTools,
     Edge               from TopoDS,
     Prism            from BRepSweep,     
     Shape           from TopoDS,
     Face            from TopoDS,
     SequenceOfCurve from TColGeom, 
     ListOfShape     from TopTools,
     Curve           from Geom, 
     Vec             from gp,
     Dir             from gp,
     Ax1             from gp,
     Plane           from Geom,     
     Pnt             from gp

raises NoSuchObject from Standard,
       NotDone      from StdFail

is

    Create 
     
    	returns  RevolutionForm  from  LocOpe;
 
    Create (Base  : Shape       from  TopoDS;
    	    Axe   : Ax1         from  gp;
	    Angle : Real        from  Standard)
	    
	returns RevolutionForm from LocOpe;     


    Perform(me:  in  out;  Base : Shape       from  TopoDS;
		    	   Axe  : Ax1         from  gp;
		           Angle: Real        from  Standard)

	is  static;


     FirstShape(me)
    
    	returns Shape from TopoDS
	---C++: return const &
	is static;


    LastShape(me)
    
    	returns Shape from TopoDS
	---C++: return const &
	is static;


    Shape(me)
    
    	returns Shape from TopoDS 
	raises  NotDone  from  StdFail
	---C++: return const &
	is static;


    Shapes(me; S: Shape from TopoDS)
    
    	returns ListOfShape from TopTools
	---C++: return const &
    	raises NoSuchObject from Standard
	       -- The exception is raised if S is not a subshape of the profile
	is static;

    IntPerf(me:  in  out) 
     
    	is  static  private;
 

fields

    myBase       : Shape             from TopoDS;
    myVec        : Vec               from gp; 
    myTra        : Vec               from gp; 
    myAngle      : Real              from Standard;
    myAxis       : Ax1               from gp;
    myAngTra     : Real              from Standard;
    myDone       : Boolean           from Standard; 
    myIsTrans    : Boolean           from Standard;     
    myRes        : Shape             from TopoDS;
    myFirstShape : Shape             from TopoDS;
    myLastShape  : Shape             from TopoDS;
    myMap        : DataMapOfShapeListOfShape    from TopTools;
    myPnt1       : Pnt               from gp;
    myPnt2       : Pnt               from gp;    
    
end RevolutionForm;     
