-- File:	RWStepFEA_RWFeaTangentialCoefficientOfLinearThermalExpansion.cdl
-- Created:	Thu Dec 12 17:51:06 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFeaTangentialCoefficientOfLinearThermalExpansion from RWStepFEA

    ---Purpose: Read & Write tool for FeaTangentialCoefficientOfLinearThermalExpansion

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FeaTangentialCoefficientOfLinearThermalExpansion from StepFEA

is
    Create returns RWFeaTangentialCoefficientOfLinearThermalExpansion from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FeaTangentialCoefficientOfLinearThermalExpansion from StepFEA);
	---Purpose: Reads FeaTangentialCoefficientOfLinearThermalExpansion

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FeaTangentialCoefficientOfLinearThermalExpansion from StepFEA);
	---Purpose: Writes FeaTangentialCoefficientOfLinearThermalExpansion

    Share (me; ent : FeaTangentialCoefficientOfLinearThermalExpansion from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFeaTangentialCoefficientOfLinearThermalExpansion;
