-- File:	GeomFill_GuideTrihedronPlan.cdl
-- Created:	Tue Jun 23 15:36:58 1998
-- Author:	Stephanie HUMEAU
--		<shu@sun17>
---Copyright:	 Matra Datavision 1998

 
class  GuideTrihedronPlan  from  GeomFill  


---Purpose: Trihedron in  the case of sweeping along a guide curve defined
-- by the orthogonal  plan on  the trajectory


inherits  TrihedronWithGuide  from  GeomFill      
    
uses  
    Shape  from  GeomAbs, 
    Array1OfReal   from TColStd, 
    HArray2OfPnt2d   from TColgp, 
    Vec  from  gp,  
    Curve  from  Geom, 
    HCurve  from  Adaptor3d, 
    TrihedronLaw  from  GeomFill, 
    Frenet  from  GeomFill,   
    PipeError  from  GeomFill,
    Vector  from  math 

raises
    OutOfRange,  ConstructionError

is 
    Create (theGuide  :  HCurve  from  Adaptor3d)   
    returns  GuideTrihedronPlan  from  GeomFill;  
     
    Init (me  :  mutable) 
    is  static  private; 
     
    SetCurve(me:mutable;  
    	     thePath  :  HCurve  from  Adaptor3d) 
    is  redefined;     
	     
    Copy(me)  returns  TrihedronLaw  from  GeomFill          
     is  redefined;
 
    ErrorStatus(me)   
    ---Purpose:Give a status to the Law              
    --         Returns PipeOk (default implementation) 
    returns  PipeError  from  GeomFill 
    is  redefined;   
        
       
    Guide(me)   
    returns  HCurve  from  Adaptor3d 
    is  redefined;      
     
    D0( me : mutable;  
        Param  : Real; 
        Tangent    : out  Vec  from  gp; 
        Normal     : out  Vec  from  gp;  
        BiNormal   : out  Vec  from  gp)        
    returns Boolean  is  redefined;    

    D1( me : mutable;  
        Param  : Real; 
        Tangent    : out  Vec  from  gp; 
    	DTangent   : out  Vec  from  gp; 
        Normal     : out  Vec  from  gp;  
        DNormal    : out  Vec  from  gp;  
        BiNormal   : out  Vec  from  gp; 
        DBiNormal  : out  Vec  from  gp)        
    returns Boolean  is  redefined;  
    
    D2( me : mutable;  
        Param  : Real; 
        Tangent    : out  Vec  from  gp; 
    	DTangent   : out  Vec  from  gp; 
    	D2Tangent  : out  Vec  from  gp; 
        Normal     : out  Vec  from  gp;  
        DNormal    : out  Vec  from  gp;  
        D2Normal   : out  Vec  from  gp;  
        BiNormal   : out  Vec  from  gp; 
        DBiNormal  : out  Vec  from  gp; 
        D2BiNormal : out  Vec  from  gp)        
    returns Boolean  is  redefined;  

       
--
--  =================== Management  of  continuity  ===================
--                 
   SetInterval(me: mutable; First, Last: Real from Standard)    
	---Purpose: Sets the bounds of the parametric interval on 
	--          the function
	--          This determines the derivatives in these values if the
	--          function is not Cn.
   is redefined;  

    NbIntervals(me; S : Shape from GeomAbs) 
	---Purpose: Returns  the number  of  intervals for  continuity
	--          <S>. 
        --          May be one if Continuity(me) >= <S>
    returns Integer  is  redefined;
 
    Intervals(me; T : in out Array1OfReal from TColStd; 
    	         S : Shape from GeomAbs)
	---Purpose: Stores in <T> the  parameters bounding the intervals
	--          of continuity <S>.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
    raises
    	OutOfRange from Standard 
    is redefined;  
  
--  ===================  To help   computation of  Tolerance   ===============	 
    GetAverageLaw(me  :  mutable;
      ATangent    : out  Vec  from  gp; 
      ANormal     : out  Vec  from  gp; 
      ABiNormal   : out  Vec  from  gp) 
     ---Purpose: Get average value of M(t) and V(t) it is usfull to 
     --          make fast approximation of rational  surfaces.        
  is  redefined;

--   =================== To help Particular case   ===============	 
    IsConstant(me) 
    ---Purpose: Say if the law is Constant

    --          Return False by Default.        
    returns  Boolean   
    is redefined;  
     
     
    IsOnlyBy3dCurve(me) 
     ---Purpose: Say if the law is defined, only by the 3d Geometry of
     --          the setted Curve  
     --          Return False by Default.        
    returns  Boolean   
    is redefined; 
     
    Origine(me  :  mutable; 
    	    OrACR1  :  Real; 
    	    OrACR2  :  Real) 
    is  redefined;
   
    InitX(me  :  mutable; 
    	  Param  :  Real  from  Standard) 
    is  private;    


fields   
    myTrimmed  :  HCurve  from  Adaptor3d;  
    myCurve  :  HCurve  from  Adaptor3d;  
    Pole  : HArray2OfPnt2d from TColgp;
    X,   XTol  :  Vector  from  math; 
    Inf,  Sup     :  Vector  from  math;
    frenet  :  Frenet  from  GeomFill;
    myNbPts  :  Integer  from  Standard;  
    myStatus  : PipeError  from  GeomFill; 
end  GuideTrihedronPlan; 
