-- File:	IGESSolid_ToolManifoldSolid.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolManifoldSolid  from IGESSolid

    ---Purpose : Tool to work on a ManifoldSolid. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses ManifoldSolid from IGESSolid,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolManifoldSolid;
    ---Purpose : Returns a ToolManifoldSolid, ready to work


    ReadOwnParams (me; ent : mutable ManifoldSolid;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : ManifoldSolid;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : ManifoldSolid;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a ManifoldSolid <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : ManifoldSolid) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : ManifoldSolid;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : ManifoldSolid; entto : mutable ManifoldSolid;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : ManifoldSolid;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolManifoldSolid;
