-- File:        Vertex.cdl
-- Created:     Fri Dec  1 11:11:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class Vertex from StepShape 

inherits TopologicalRepresentationItem from StepShape 

uses

	HAsciiString from TCollection
is

	Create returns mutable Vertex;
	---Purpose: Returns a Vertex


end Vertex;
