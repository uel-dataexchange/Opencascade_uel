-- File:        SurfaceModel.cdl
-- Created:     Fri Dec  1 11:11:11 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class SurfaceModel from StepShape inherits SelectType from StepData

	-- <SurfaceModel> is an EXPRESS Select Type construct translation.
	-- it gathers : ShellBasedSurfaceModel, FaceBasedSurfaceModel
	-- Rev4 : only remains ShellBasedSurfaceModel

uses

	ShellBasedSurfaceModel
--	FaceBasedSurfaceModel
is

	Create returns SurfaceModel;
	---Purpose : Returns a SurfaceModel SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a SurfaceModel Kind Entity that is :
	--        1 -> ShellBasedSurfaceModel
	--        2 -> FaceBasedSurfaceModel
	--        0 else

	ShellBasedSurfaceModel (me) returns any ShellBasedSurfaceModel;
	---Purpose : returns Value as a ShellBasedSurfaceModel (Null if another type)

end SurfaceModel;

