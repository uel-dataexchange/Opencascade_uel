-- File:	StepWriter.cdl
-- Created:	Tue Feb 11 19:54:04 1992
-- Author:	Christian CAILLET
--		<cky@phobox>
---Copyright:	 Matra Datavision 1992


class StepWriter  from StepData

    ---Purpose : manages atomic file writing, under control of StepModel (for
    --           general organisation of file) and each class of Transient
    --           (for its own parameters) : prepares text to be written then
    --           writes it
    --           A stream cannot be used because Step limits line length at 72
    --           In more, a specific object offers more appropriate functions

uses Integer, Boolean, Real, Character, Transient, Logical from StepData,     -- OStream,
     AsciiString from TCollection,  HAsciiString from TCollection,
     HSequenceOfHAsciiString,  HArray1OfInteger,
     LineBuffer, FloatWriter, CheckIterator,
     StepModel, WriterLib, Protocol from StepData,
     SelectMember from StepData, Field from StepData, PDescr from StepData,
     FieldList from StepData, ESDescr from StepData,
     HArray1OfReal from TColStd

raises InterfaceMismatch

is

    Create (amodel : StepModel) returns StepWriter;
    ---Purpose : Creates an empty StepWriter from a StepModel. The StepModel
    --           provides the Number of Entities, as identifiers for File

    	--  Options for Sending Forms  --

    LabelMode (me : in out) returns Integer;
    ---Purpose : ModeLabel controls how to display entity ids :
    --           0 (D) gives entity number in the model
    --           1 gives the already recorded label (else, its number)
    --  Warning : conflicts are not controlled
    ---C++ : return &

    TypeMode  (me : in out) returns Integer;
    ---Purpose : TypeMode  controls the type form to use :
    --           0 (D) for normal long form
    --           1 for short form (if a type name has no short form, normal
    --             long form is then used)
    ---C++ : return &

    FloatWriter (me : in out) returns FloatWriter;
    ---Purpose : Returns the embedded FloatWriter, which controls sending Reals
    --           Use this method to access FloatWriter in order to consult or
    --           change its options (MainFormat, FormatForRange,ZeroSuppress),
    --           because it is returned as the address of its field
    ---C++ : return &

    	-- --  Description of Scopes  -- --   (to be done before sending)

    SetScope (me : in out; numscope,numin : Integer)
    ---Purpose : Declares the Entity Number <numscope> to correspond to a Scope
    --           which contains the Entity Number <numin>. Several calls to the
    --           same <numscope> add Entities in this Scope, in this order.
    	raises InterfaceMismatch;
    ---Purpose:           Error if <numin> is already declared in the Scope
    --  Warning : the declaration of the Scopes is assumed to be consistent,
    --           i.e. <numin> is not referenced from outside this Scope
    --           (not checked here)

    IsInScope (me; num : Integer) returns Boolean;
    ---Purpose : Returns True if an Entity identified by its Number is in a Scope

    	-- --  Sending Parts of a Model  -- --

    SendModel  (me : in out; protocol : Protocol from StepData;
    	    	    	     headeronly : Boolean = Standard_False)
    ---Purpose : Sends the complete Model, included HEADER and DATA Sections
    --           Works with a WriterLib defined through a Protocol
    --           If <headeronly> is given True, only the HEADER Section is sent
    --           (used to Dump the Header of a StepModel)
      raises InterfaceMismatch;
    --           Error if any of the called Send's falls in Error

    SendHeader (me : in out);
    ---Purpose : Begins model header

    SendData (me : in out) raises InterfaceMismatch;
    ---Purpose : Begins data section; error if EndSec was not set

    SendEntity (me : in out; nument : Integer; lib : WriterLib)
    ---Purpose : Send an Entity of the Data Section. If it corresponds to a
    --           Scope, also Sends the Scope informations and contained Items
      raises InterfaceMismatch;
    --           Error if any of the called Send's falls in Error

    EndSec (me : in out);
    ---Purpose : sets end of section; to be done before passing to next one

    EndFile (me : in out)  raises InterfaceMismatch;
    ---Purpose : sets end of file; error is EndSec was not set

    	-- --   Managing line   -- --

    AddString (me : in out; str : AsciiString from TCollection; more : Integer = 0)
    	is private;
    ---Purpose : adds a string to current line; first flushes it if full
    --           (72 char); more allows to ask a reserve at end of line : flush
    --           is done if remaining length (to 72) is less than <more>

    AddString (me : in out; str : CString; lnstr : Integer; more : Integer = 0)
    	is private;
    ---Purpose : Same as above, but the string is given by CString + Length


    NewLine (me : in out; evenempty : Boolean);
    ---Purpose : flushes current line; if empty, flushes it (defines a new
    --           empty line) if evenempty is True; else, skips it

    JoinLast (me : in out; newline : Boolean);
    ---Purpose : joins current line to last one, only if new length is 72 max
    --           if newline is True, a new current line begins; else, current
    --           line is set to the last line (once joined) itself an can be
    --           completed

    Indent (me : in out; onent : Boolean);
    ---Purpose : asks that further indentations will begin at position of
    --           entity first opening bracket; else they begin at zero (def)
    --           for each sublist level, two more blancks are added at beginning
    --           (except for text continuation, which must begin at true zero)

    	-- --   Sending entities   -- --

    SendIdent (me : in out; ident : Integer);
    ---Purpose : begins an entity with an ident plus '=' (at beginning of line)
    --           entity ident is its Number given by the containing Model
    --  Warning : <ident> must be, either Number or Label, according LabelMode

    SendScope (me : in out);
    ---Purpose : sets a begin of Scope (ends this line)

    SendEndscope (me : in out);
    ---Purpose : sets an end of Scope  (on a separate line)

    Comment (me : in out; mode : Boolean);
    ---Purpose : sets a comment mark : if mode is True, begins Comment zone,
    --           if mode is False, ends Comment zone (if one is begun)

    SendComment (me : in out; text : HAsciiString from TCollection)
      raises InterfaceMismatch;
    ---Purpose : sends a comment. Error if we are not inside a comment zone

    SendComment (me : in out; text : CString)  raises InterfaceMismatch;
    ---Purpose : same as above but accepts a CString (ex.: "..." directly)

    StartEntity (me : in out; atype : AsciiString from TCollection);
    ---Purpose : sets entity's StepType, opens brakets, starts param no to 0
    --           params are separated by comma
    --           Remark : for a Multiple Type Entity (see Express ANDOR clause)
    --           StartComplex must be called before sending componants, then
    --           each "Componant" must be send separately (one call to
    --           StartEntity for each one) : the Type which preceeds is then
    --           automaticaly closed. Once all the componants have been sent,
    --           EndComplex must be called, then and only then EndEntity

    StartComplex (me : in out);
    ---Purpose : sends the start of a complex entity, which is a simple open
    --           bracket (without increasing braket level)
    --           It must be called JUST AFTER SendEntity and BEFORE sending
    --           componants, each one begins by StartEntity

    EndComplex   (me : in out);
    ---Purpose : sends the end of a complex entity : a simple closed bracket
    --           It must be called AFTER sending all the componants and BEFORE
    --           the final call to EndEntity

    	-- --   Sending Parameters   -- --

    SendField  (me : in out; fild : Field; descr : PDescr);
    ---Purpose : Sends the content of a field, controlled by its descriptor
    --           If the descriptor is not defined, follows the description
    --           detained by the field itself

    SendSelect (me : in out; sm : SelectMember; descr : PDescr);
    ---Purpose : Sends a SelectMember, which cab be named or not

    SendList   (me : in out; list : FieldList; descr : ESDescr);
    ---Purpose : Send the content of an entity as being a FieldList controlled
    --           by its descriptor. This includes start and end brackets but
    --           not the entity type

    OpenSub (me : in out);
    ---Purpose : open a sublist by a '('

    OpenTypedSub (me : in out; subtype : CString);
    ---Purpose : open a sublist with its type then a '('

    CloseSub (me : in out);
    ---Purpose : closes a sublist by a ')'

    AddParam (me : in out);
    ---Purpose : prepares adding a parameter (that is, adds ',' except for
    --           first one); normally for internal use; can be used to send
    --           a totally empty parameter (with no litteral value)

    Send (me : in out; val : Integer);
    ---Purpose : sends an integer parameter

    Send (me : in out; val : Real);
    ---Purpose : sends a real parameter (wroks with FloatWriter)

    Send (me : in out; val : AsciiString from TCollection);
    ---Purpose : sends a text given as string (it will be set between '...')

    Send (me : in out; val : Transient);
    ---Purpose : sends a reference to an entity (its identifier with '#')
    --           REMARK 1 : a Null <val> is interpreted as "Undefined"
    --           REMARK 2 : for an HAsciiString which is not recorded in the
    --           Model, it is send as its String Content, between quotes

    SendBoolean (me : in out; val : Boolean);
    ---Purpose : sends a Boolean as .T. for True or .F. for False
    --           (it is an useful case of Enum, which is built-in)

    SendLogical (me : in out; val : Logical from StepData);
    ---Purpose : sends a Logical as .T. or .F. or .U. according its Value
    --           (it is a standard case of Enum for Step, and is built-in)

    SendString (me : in out; val : AsciiString from TCollection);
    ---Purpose : sends a string exactly as it is given

    SendString (me : in out; val : CString);
    ---Purpose : sends a string exactly as it is given

    SendEnum (me : in out; val : AsciiString from TCollection);
    ---Purpose : sends an enum given by String (litteral expression)
    --           adds '.' around it if not done
    --           Remark : val can be computed by class EnumTool from StepData:
    --             StepWriter.SendEnum (myenum.Text(enumval));

    SendEnum (me : in out; val : CString);
    ---Purpose : sends an enum given by String (litteral expression)
    --           adds '.' around it if not done

    SendArrReal(me : in out; anArr : HArray1OfReal from TColStd);
    ---Purpose : sends an array of real

    SendUndef (me : in out);
    ---Purpose : sends an undefined (optionnal absent) parameter (by '$')

    SendDerived (me : in out);
    ---Purpose : sends a "Derived" parameter (by '*'). A Derived Parameter has
    --           been inherited from a Super-Type then redefined as being
    --           computed by a function. Hence its value in file is senseless.

    EndEntity (me : in out) raises InterfaceMismatch;
    ---Purpose : sends end of entity (closing bracket plus ';')
    --           Error if count of opened-closed brackets is not null

    	-- --   Printing on an output   -- --

    CheckList (me) returns CheckIterator;
    ---Purpose : Returns the check-list, which has received possible checks :
    --           for unknown entities, badly loaded ones, null or unknown
    --           references

    NbLines (me) returns Integer;
    ---Purpose : Returns count of Lines

    Line (me; num : Integer) returns HAsciiString from TCollection;
    ---Purpose : Returns a Line given its rank in the File

    Print (me : in out; S : in out OStream) returns Boolean;
    ---Purpose : writes result on an output defined as an OStream
    --           then clears it

fields

    themodel  : StepModel;
    thefile   : HSequenceOfHAsciiString;
    thecurr   : LineBuffer;
    thesect   : Boolean;  -- False at very start or after EndSec
    thecomm   : Boolean;  -- are we in inside a comment
    thefirst  : Boolean;  -- True on first parameter, False on following ones
    themult   : Boolean;  -- True after sending first type (for Multiple Type)
    thelevel  : Integer;  -- current sublist level
    theindent : Boolean;  -- True to indent at entity opening bracket
    theindval : Integer;  -- position of entity opening bracket

    thetypmode   : Integer;
    thefloatw : FloatWriter;  -- control of sending Reals

    thechecks    : CheckIterator;
    thenum       : Integer;

    thelabmode   : Integer;
    thescopebeg  : HArray1OfInteger;
    thescopeend  : HArray1OfInteger;
    thescopenext : HArray1OfInteger;

end StepWriter;
