-- File:	RWStepAP214_RWClass.cdl
-- Created:	Wed May 10 15:09:06 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWClass from RWStepAP214

    ---Purpose: Read & Write tool for Class

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    Class from StepAP214

is
    Create returns RWClass from RWStepAP214;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : Class from StepAP214);
	---Purpose: Reads Class

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: Class from StepAP214);
	---Purpose: Writes Class

    Share (me; ent : Class from StepAP214;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWClass;
