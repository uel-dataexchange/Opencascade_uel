-- File:	TopOpeBRepTool_PurgeInternalEdges.cdl
-- Created:	Thu Nov 19 15:23:38 1998
-- Author:	Jean-Michel BOULCOURT
--		<jmb@coulox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1998


class PurgeInternalEdges from TopOpeBRepTool 

	---Purpose: remove from  a shape, the  internal edges that are
	--          not  connected to any face in  the shape.   We can
	--             get  the    list   of      the    edges  as   a
	--          DataMapOfShapeListOfShape with a Face of the Shape
	--          as  the key and  a  list of internal  edges as the
	--           value.  The list   of internal edges  means edges
	--          that are  not connected to any  face in the shape.
	--          
	--          Example of use          :
	--               TopTools_DataMapOfShapeListOfShape     mymap;
	--               TopOpeBRepTool_PurgeInternalEdges
	--               mypurgealgo(mysolid); mypurgealgo.GetFaces(mymap);
	--            

uses
  Shape from TopoDS,
  DataMapOfShapeListOfShape from TopTools,
  IndexedDataMapOfShapeListOfShape from TopTools
  
  raises
      	ConstructionError from Standard,
        NullObject        from Standard

is

    Create (theShape : Shape from TopoDS;
    	    PerformNow : Boolean from Standard = Standard_True)
    returns PurgeInternalEdges from TopOpeBRepTool
    raises NullObject        from Standard, 
           ConstructionError from Standard;
        ---Purpose: Initialize   members and  begin  exploration   of  shape
        --          depending of the value of PerformNow

    Faces (me : in out ; theMapFacLstEdg : in out DataMapOfShapeListOfShape from TopTools);
    	---Purpose: returns  the list  internal edges associated  with
    	--          the faces of the  myShape. If PerformNow was False
    	--          when created, then call the private Perform method
    	--          that do the main job.

    Shape (me : in out)
    returns Shape from TopoDS
    raises NullObject        from Standard;
    	---Purpose: returns myShape modified with the list of internal
    	--          edges removed from it.
        ---C++: return &
    
    NbEdges (me )
    returns Integer from Standard
    raises NullObject        from Standard;
    	---Purpose: returns the number of edges candidate to be removed
    	---C++: return const


    IsDone (me)  
    returns Boolean from Standard
        ---Purpose: returns False  if the list  of internal  edges has
        --          not been extracted
        ---C++: inline
    is static;
    
    Perform (me : in out);
    ---Purpose:  Using   the list  of internal edge    from each face,
    --           rebuild myShape by removing thoses edges.
    --          

    BuildList (me : in out)
    ---Purpose: Do the main job. Explore all the  edges of myShape and
    --          build a map with  faces as a key  and list of internal
    --          edges(without connected faces) as value.
    --          
    is private;

fields

  myShape         : Shape from TopoDS;
  myIsDone        : Boolean from Standard;
  myMapFacLstEdg  : DataMapOfShapeListOfShape from TopTools;
  myMapEdgLstFac  : IndexedDataMapOfShapeListOfShape from TopTools is protected;
  
end PurgeInternalEdges;
