-- File:	StepRepr_ConfigurationDesignItem.cdl
-- Created:	Fri Nov 26 16:26:26 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class ConfigurationDesignItem from StepRepr
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type ConfigurationDesignItem

uses
    ProductDefinition from StepBasic,
    ProductDefinitionFormation from StepBasic

is
    Create returns ConfigurationDesignItem from StepRepr;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of ConfigurationDesignItem select type
	--          1 -> ProductDefinition from StepBasic
	--          2 -> ProductDefinitionFormation from StepBasic
	--          0 else

    ProductDefinition (me) returns ProductDefinition from StepBasic;
	---Purpose: Returns Value as ProductDefinition (or Null if another type)

    ProductDefinitionFormation (me) returns ProductDefinitionFormation from StepBasic;
	---Purpose: Returns Value as ProductDefinitionFormation (or Null if another type)

end ConfigurationDesignItem;
