-- File:	StepShape_NonManifoldSurfaceShapeRepresentation.cdl
-- Created:	Fri Dec 28 16:02:02 2001 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class NonManifoldSurfaceShapeRepresentation from StepShape
inherits ShapeRepresentation from StepShape

    ---Purpose: Representation of STEP entity NonManifoldSurfaceShapeRepresentation

uses
    HAsciiString from TCollection,
    HArray1OfRepresentationItem from StepRepr,
    RepresentationContext from StepRepr

is
    Create returns NonManifoldSurfaceShapeRepresentation from StepShape;
	---Purpose: Empty constructor

end NonManifoldSurfaceShapeRepresentation;
