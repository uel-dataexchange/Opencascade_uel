-- File:	StepToGeom.cdl
-- Created:	Fri Jun 11 18:17:21 1993
-- Author:	Martine LANGLOIS
---Copyright:	 Matra Datavision 1993

package StepToGeom

--- Purpose: Creation des entites geometriques de Geom a partir du schema 
--  StepGeom (Part42, geometric)

uses  gp, Geom, Geom2d, StepGeom, StdFail

is

private deferred class Root;
class MakeCartesianPoint;
class MakeCartesianPoint2d;
class MakeAxisPlacement;
class MakeAxis1Placement;
class MakeAxis2Placement;
class MakeDirection;
class MakeDirection2d;
class MakeVectorWithMagnitude;
class MakeVectorWithMagnitude2d;
class MakeCurve;
class MakeTrimmedCurve;
class MakeTrimmedCurve2d;
class MakeCurve2d;
class MakeConic;
class MakeConic2d;
class MakeBoundedCurve;
class MakeBoundedCurve2d;
class MakeEllipse;
class MakeEllipse2d;
class MakeHyperbola;
class MakeHyperbola2d;
class MakeParabola;
class MakeParabola2d;
class MakeCircle;
class MakeCircle2d;
class MakeBSplineCurve;
class MakeBSplineCurve2d;
class MakeLine;
class MakeLine2d;
class MakePolyline;
class MakePolyline2d;
class MakePlane;
class MakeSurface;
class MakeBoundedSurface;
class MakeElementarySurface;
class MakeSweptSurface;
class MakeConicalSurface;
class MakeCylindricalSurface;
class MakeRectangularTrimmedSurface;
class MakeSphericalSurface;
class MakeSurfaceOfLinearExtrusion;
class MakeSurfaceOfRevolution;
class MakeToroidalSurface;
class MakeBSplineSurface;
class MakeTransformation3d;
class MakeTransformation2d;

-- class CheckSurfaceClosure;

end StepToGeom;
