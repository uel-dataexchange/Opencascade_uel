-- File:	MDocStd_XLinkRetrievalDriver.cdl
--      	-----------------------------
-- Author:	DAUTRY Philippe
--		<fid@fox.paris1.matra-dtv.fr>
---Copyright:	 MATRA DATAVISION 1997

---Version:	0.0
---History:	Version	Date		Purpose
--		0.0	Sep 17 1997	Creation


class XLinkRetrievalDriver from MDocStd
    inherits ARDriver from MDF

	---Purpose: Tool used to translate a persistent XLink into a
	--          transient one.

uses

    RRelocationTable from MDF,
    Attribute        from TDF,
    Attribute        from PDF, 
    MessageDriver    from CDM

is

    Create (theMessageDriver : MessageDriver from CDM) -- Version 0
    returns mutable XLinkRetrievalDriver from MDocStd;

    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type XLink from PXref.

    NewEmpty (me)
    returns mutable Attribute from TDF;


    Paste(me;
    	  aSource     :          Attribute        from PDF;
    	  aTarget     : mutable  Attribute        from TDF;
    	  aRelocTable :          RRelocationTable from MDF);


end XLinkRetrievalDriver from MDocStd;
