-- File:        AutoDesignDateAndPersonItem.cdl
-- Created:     Fri Dec  1 11:11:10 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class AutoDesignDateAndPersonItem from StepAP214 inherits SelectType from StepData

	-- <AutoDesignDateAndPersonItem> is an EXPRESS Select Type construct translation.
	-- it gathers : Product, ProductDefinition, ProductDefinitionFormation, Representation
	-- Rev4 adds : AutoDesignOrganizationAssignment


uses
     AutoDesignOrganizationAssignment from StepAP214,
     Product from StepBasic,
     ProductDefinition from StepBasic,
     ProductDefinitionFormation from StepBasic,
     Representation from StepRepr,
     AutoDesignDocumentReference from StepAP214,
     ExternallyDefinedRepresentation from StepRepr,
     ProductDefinitionRelationship from StepBasic,
     ProductDefinitionWithAssociatedDocuments from StepBasic

is

	Create returns AutoDesignDateAndPersonItem;
	---Purpose : Returns a AutoDesignDateAndPersonItem SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a AutoDesignDateAndPersonItem Kind Entity that is :
	-- 1     AutoDesignOrganizationAssignment from StepAP214,
	-- 2     Product from StepBasic,
	-- 3     ProductDefinition from StepBasic,
	-- 4     ProductDefinitionFormation from StepBasic,
	-- 5     Representation from StepRepr,
	-- 6     AutoDesignDocumentReference from StepAP214,
	-- 7     ExternallyDefinedRepresentation from StepRepr,
	-- 8     ProductDefinitionRelationship from StepBasic,
	-- 9     ProductDefinitionWithAssociatedDocuments from StepBasic
	--        0 else

     AutoDesignOrganizationAssignment (me) returns AutoDesignOrganizationAssignment from StepAP214;
     Product (me) returns Product from StepBasic;
     ProductDefinition (me) returns ProductDefinition from StepBasic;
     ProductDefinitionFormation (me) returns ProductDefinitionFormation from StepBasic;
     Representation (me) returns Representation from StepRepr;
     AutoDesignDocumentReference (me) returns AutoDesignDocumentReference from StepAP214;
     ExternallyDefinedRepresentation (me) returns ExternallyDefinedRepresentation from StepRepr;
     ProductDefinitionRelationship (me) returns ProductDefinitionRelationship from StepBasic;
     ProductDefinitionWithAssociatedDocuments (me) returns ProductDefinitionWithAssociatedDocuments from StepBasic;

end AutoDesignDateAndPersonItem;

