-- File:        UniformCurve.cdl
-- Created:     Fri Dec  1 11:11:30 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class UniformCurve from StepGeom 

inherits BSplineCurve from StepGeom 

uses

	HAsciiString from TCollection, 
	Integer from Standard, 
	HArray1OfCartesianPoint from StepGeom, 
	BSplineCurveForm from StepGeom, 
	Logical from StepData
is

	Create returns mutable UniformCurve;
	---Purpose: Returns a UniformCurve


end UniformCurve;
