-- File:	BRepTools_TrsfModification.cdl
-- Created:	Thu Aug 25 16:38:07 1994
-- Author:	Jacques GOUSSARD
--		<jag@ecolox>
---Copyright:	 Matra Datavision 1994


class TrsfModification from BRepTools inherits Modification from BRepTools

---Purpose: Describes a modification that uses a gp_Trsf to
-- change the geometry of a shape. All functions return
-- true and transform the geometry of the shape.
        
uses Face     from TopoDS,
     Edge     from TopoDS,
     Vertex   from TopoDS,
     Location from TopLoc,
     Shape    from GeomAbs,
     
     Surface  from Geom,
     Curve    from Geom,
     Curve    from Geom2d,
     
     Trsf     from gp,
     Pnt      from gp
     
is

    Create (T : Trsf from gp) returns mutable TrsfModification from BRepTools; 
    
    Trsf(me: mutable)
	---Purpose: Provides access to the gp_Trsf associated with this
    	-- modification. The transformation can be changed.
    		---C++: return &
    	returns Trsf from gp
	is static;


    NewSurface(me: mutable; F       :     Face     from TopoDS;
                            S       : out Surface  from Geom;
		            L       : out Location from TopLoc;
		            Tol     : out Real     from Standard;
                            RevWires : out Boolean from Standard;
                            RevFace  : out Boolean from Standard)
    
      	---Purpose: Returns true if the face F has been modified.
-- If the face has been modified:
-- - S is the new geometry of the face,
-- - L is its new location, and
-- - Tol is the new tolerance.
-- RevWires is set to true when the modification
-- reverses the normal of the surface (the wires have to be reversed).
-- RevFace is set to true if the orientation of the
-- modified face changes in the shells which contain it.
-- For this class, RevFace returns true if the gp_Trsf
-- associated with this modification is negative.
    
    
    	returns Boolean from Standard
	;
	

    NewCurve(me: mutable; E  :     Edge     from TopoDS;
                          C  : out Curve    from Geom;
		          L  : out Location from TopLoc;
		          Tol: out Real     from Standard)
    
    	returns Boolean from Standard
	;
	
	---Purpose: Returns true if the edge E has been modified.
-- If the edge has been modified:
-- - C is the new geometric support of the edge,
-- - L is the new location, and
-- - Tol is the new tolerance.
--   If the edge has not been modified, this function
-- returns false, and the values of C, L and Tol are not significant.
    

    NewPoint(me: mutable; V  :     Vertex   from TopoDS;
                          P  : out Pnt      from gp;
		          Tol: out Real     from Standard)
    
    	returns Boolean from Standard
	;
	
	---Purpose: Returns true if the vertex V has been modified.
-- If the vertex has been modified:
-- - P is the new geometry of the vertex, and
-- - Tol is the new tolerance.
--   If the vertex has not been modified this function
-- returns false, and the values of P and Tol are not significant.
    

    NewCurve2d(me: mutable;  E    :     Edge     from TopoDS;
                             F    :     Face     from TopoDS;
                             NewE :     Edge     from TopoDS;
                             NewF :     Face     from TopoDS;
                             C    : out Curve    from Geom2d;
		             Tol  : out Real     from Standard)
    
    	returns Boolean from Standard
	;
	
	---Purpose: Returns true if the edge E has a new curve on surface on the face F.
-- If a new curve exists:
-- - C is the new geometric support of the edge,
-- - L is the new location, and
-- - Tol the new tolerance.
--   If no new curve exists, this function returns false, and
-- the values of C, L and Tol are not significant.
    

    NewParameter(me: mutable; V  :     Vertex   from TopoDS;
                              E  :     Edge     from TopoDS;
                              P  : out Real     from Standard;
  		              Tol: out Real     from Standard)
    
    	returns Boolean from Standard
	;
	
	---Purpose: Returns true if the Vertex V has a new parameter on the edge E.
-- If a new parameter exists:
-- - P is the parameter, and
-- - Tol is the new tolerance.
--   If no new parameter exists, this function returns false,
-- and the values of P and Tol are not significant.
    


    

    Continuity(me: mutable; E          : Edge from TopoDS;
    	                    F1,F2      : Face from TopoDS;
			    NewE       : Edge from TopoDS;
			    NewF1,NewF2: Face from TopoDS)
    
    	returns Shape from GeomAbs
	
	---Purpose: Returns the  continuity of  <NewE> between <NewF1>
	--          and <NewF2>.
	--          
	--          <NewE> is the new  edge created from <E>.  <NewF1>
	--          (resp. <NewF2>) is the new  face created from <F1>
	--          (resp. <F2>).

    	;



fields

    myTrsf : Trsf from gp;

end TrsfModification;
