-- File:	IGESSolid_ToolEllipsoid.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolEllipsoid  from IGESSolid

    ---Purpose : Tool to work on a Ellipsoid. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses Ellipsoid from IGESSolid,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolEllipsoid;
    ---Purpose : Returns a ToolEllipsoid, ready to work


    ReadOwnParams (me; ent : mutable Ellipsoid;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : Ellipsoid;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : Ellipsoid;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a Ellipsoid <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : Ellipsoid) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : Ellipsoid;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : Ellipsoid; entto : mutable Ellipsoid;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : Ellipsoid;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolEllipsoid;
