-- File:	StepBasic_DocumentUsageConstraint.cdl
-- Created:	Tue Jun 30 15:07:15 1998
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1998


class DocumentUsageConstraint  from StepBasic    inherits TShared from MMgt

uses
     Document from StepBasic,
     HAsciiString from TCollection

is

    Create returns mutable DocumentUsageConstraint;

    Init (me : mutable;
    	  aSource : Document;
	  ase  : HAsciiString;
	  asev : HAsciiString);

    Source (me) returns Document;
    SetSource (me : mutable; aSource : Document);

    SubjectElement (me) returns HAsciiString;
    SetSubjectElement (me : mutable; ase : HAsciiString);

    SubjectElementValue (me) returns HAsciiString;
    SetSubjectElementValue (me : mutable; asev : HAsciiString);

fields

    theSource : Document;
    theSE  : HAsciiString;
    theSEV : HAsciiString;

end DocumentUsageConstraint;
