-- File:	RWStepBasic_RWSiUnitAndAreaUnit.cdl
-- Created:	Mon Oct 11 15:33:17 1999
-- Author:	data exchange team
--		<det@friendox>
---Copyright:	 Matra Datavision 1999


class RWSiUnitAndAreaUnit from RWStepBasic 

	---Purpose: Read & Write Module for SiUnitAndAreaUnit

uses

    Check from Interface,
    StepReaderData from StepData,
    StepWriter from StepData,
    SiUnitAndAreaUnit from StepBasic

is

    Create returns  RWSiUnitAndAreaUnit from RWStepBasic;
    
    ReadStep (me; data: StepReaderData; num: Integer;
	          ach : in out Check;   ent: mutable SiUnitAndAreaUnit from StepBasic);
    
    WriteStep (me; SW : in out StepWriter; ent: SiUnitAndAreaUnit from StepBasic);


end RWSiUnitAndAreaUnit;
