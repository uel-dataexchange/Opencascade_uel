-- File:        Edge.cdl
-- Created:     Mon Dec  4 12:02:26 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWEdge from RWStepShape

	---Purpose : Read & Write Module for Edge

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Edge from StepShape,
     EntityIterator from Interface

is

	Create returns RWEdge;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Edge from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : Edge from StepShape);

	Share(me; ent : Edge from StepShape; iter : in out EntityIterator);

end RWEdge;
