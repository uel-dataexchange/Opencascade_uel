-- File:        QuasiUniformSurfaceAndRationalBSplineSurface.cdl
-- Created:     Mon Dec  4 12:02:34 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWQuasiUniformSurfaceAndRationalBSplineSurface from RWStepGeom

	---Purpose : Read & Write Module for QuasiUniformSurfaceAndRationalBSplineSurface

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     QuasiUniformSurfaceAndRationalBSplineSurface from StepGeom,
     EntityIterator from Interface

is

	Create returns RWQuasiUniformSurfaceAndRationalBSplineSurface;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable QuasiUniformSurfaceAndRationalBSplineSurface from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : QuasiUniformSurfaceAndRationalBSplineSurface from StepGeom);

	Share(me; ent : QuasiUniformSurfaceAndRationalBSplineSurface from StepGeom; iter : in out EntityIterator);

end RWQuasiUniformSurfaceAndRationalBSplineSurface;
