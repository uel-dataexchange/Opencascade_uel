-- File:	RWStepElement_RWCurveElementEndReleasePacket.cdl
-- Created:	Thu Dec 12 17:29:00 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWCurveElementEndReleasePacket from RWStepElement

    ---Purpose: Read & Write tool for CurveElementEndReleasePacket

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    CurveElementEndReleasePacket from StepElement

is
    Create returns RWCurveElementEndReleasePacket from RWStepElement;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : CurveElementEndReleasePacket from StepElement);
	---Purpose: Reads CurveElementEndReleasePacket

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: CurveElementEndReleasePacket from StepElement);
	---Purpose: Writes CurveElementEndReleasePacket

    Share (me; ent : CurveElementEndReleasePacket from StepElement;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWCurveElementEndReleasePacket;
