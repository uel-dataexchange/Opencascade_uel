-- File     : Prs2d.cdl
-- Created  : February  2000
-- Author   : Tanya COOL
---Copyright: Matra Datavision 2000

package Prs2d
 
 ---Purpose: package provides the graphic attribute manager Drawer,
 --          the set of aspect classes for storing hte session attributes 
 --          and default attributes for the objects. 

uses

	Graphic2d,
	Aspect,
  	Quantity,
	TShort,
	Standard,
	gp,
	Geom2d,
	TCollection,
	TColgp,
	TColStd,
	TopoDS,
	GCPnts
is
    enumeration AspectName is

        AN_UNKNOWN,
        AN_LINE,
        AN_HIDDENLINE,
        AN_TEXT,
        AN_HIDINGPOLY,
	    AN_HIDINGTEXT,
	    AN_FRAMEDTEXT,
        
    -- For new aspect types
        AN_LAST

    end AspectName;

    enumeration TypeOf2DObject is

		 TOO_UNKNOWN,
		 TOO_ANGLE,
		 TOO_ARROW,
		 TOO_CURVE,
		 TOO_DATUM,
		 TOO_DIAMETER,
		 TOO_ELLIPSERADIUS,
		 TOO_EQUALDISTANCE,
		 TOO_LENGTH
							
	end TypeOf2DObject;
			  
    enumeration ArrowSide is 

        AS_NONE, 
        AS_FIRSTAR, 
        AS_LASTAR, 
        AS_BOTHAR, 
        AS_FIRSTPT, 
        AS_LASTPT, 
        AS_BOTHPT,
        AS_FIRSTAR_LASTPT, 
        AS_FIRSTPT_LASTAR
				
	end ArrowSide;
              
    enumeration TypeOfArrow is 

        TOA_OPENED,
        TOA_CLOSED,
        TOA_FILLED
	
    end TypeOfArrow;

    enumeration TypeOfDist is 
      
	  TOD_AUTOMATIC,
	  TOD_OBLIQUE,
	  TOD_HORIZONTAL,
	  TOD_VERTICAL
	  
    end TypeOfDist;

    enumeration TypeOfAxis is 
    
	  TOAX_Unknown,
	  TOAX_XAxis,
	  TOAX_YAxis

    end TypeOfAxis;

	enumeration TypeOfTolerance is 
	   
	   TOT_TAPER,
	   TOT_SYMTOTAL,
       TOT_SYMCIRCULAR,
       TOT_SYMMETRY,
       TOT_CONCENTRIC,
	   TOT_POSITION,
       TOT_ANGULARITY,
	   TOT_PERPENDIC,
	   TOT_PARALLELISM,
	   TOT_SURFACEPROF,
	   TOT_LINEPROF,
	   TOT_CYLINDRIC,
	   TOT_CIRCULARITY,
	   TOT_FLATNESS,
	   TOT_STRAIGHTNESS,
	   TOT_NONE

	end TypeOfTolerance;
    
    enumeration TypeOfSymbol is 
      
	  TOS_NONE,
	  TOS_DIAMETER,


      TOS_LAST
	  
    end TypeOfSymbol;

    enumeration TypeOfRadius is 
      
	  TOR_STANDARD,
	  TOR_CENTER,
	  TOR_REVARROW,
	  TOR_CENTREV, 
      TOR_NONE
	  
    end TypeOfRadius;

    exception SymbolDefinitionError inherits OutOfRange;
        
    deferred class AspectRoot;
    
    -- Standard aspects

    class AspectLine;
    class AspectText;

    class AspectHidingPoly; 
    class AspectHidingText;
    class AspectFramedText;
	
	-- Standard primitives
	
	class Point;
	class Axis;
	class Arrow;

	-- Dimensions 

    deferred class Dimension;
	class Angle;
	class Length;
    class Radius;
	class Diameter;
	class Repere;
    
    class RadiusIndep;

	class ToleranceFrame;

	deferred class Tolerance;

	class Straightness;
	class Flatness;
	class Circularity;
    class Cylindric;
	class LineProfile;
	class SurfProfile;
	class Parallelism;
    class Perpendicular;
	class Angularity;
	class Position;
	class Concentric;
	class Symmetry;
	class SymTotal;
    class SymCircular;
	class Taper;

    class DrawSymbol;

    class Drawer;
 			
    class DataMapOfAspectRoot instantiates DataMap from TCollection
          ( Integer from Standard,
            AspectRoot from Prs2d,
            MapIntegerHasher from  TColStd );

end Prs2d;
