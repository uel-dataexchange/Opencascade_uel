-- File:	BezierCurve2d.cdl
-- Created:	Fri May 22 10:45:54 1992
-- Author:	Jean Claude VAUTHIER
--		<jcv@sdsun4>
---Copyright:	 Matra Datavision 1992



class BezierCurve2d


from DrawTrSurf


inherits Curve2d from DrawTrSurf


uses BezierCurve from Geom2d,
     Color from Draw,
     Display from Draw,
     Drawable3D from Draw


is


  Create (C : BezierCurve from Geom2d)
        --- Purpose :
        --  creates a drawable Bezier curve from a Bezier curve of 
        --  package Geom2d.
     returns mutable BezierCurve2d from DrawTrSurf;


  Create (C : BezierCurve from Geom2d;
          CurvColor, PolesColor : Color from Draw;
          ShowPoles : Boolean; Discret : Integer)
     returns mutable BezierCurve2d from DrawTrSurf;


  DrawOn (me; dis : in out Display from Draw)
     is redefined static;


  ShowPoles (me : mutable)
     is static;


  ClearPoles (me : mutable)
     is static;
     
  
  FindPole(me; X,Y : Real; D : Display from Draw; Prec : Real; 
           Index : in out Integer)
        --- Purpose :
        --  Returns in <Index> the index of the first pole  of the
        --  curve projected by the Display <D> at a distance lower
        --  than <Prec> from <X,Y>. If no pole  is found  index is
        --  set to 0, else index is always  greater than the input
        --  value of index.
  is static;
  
  
  SetPolesColor (me : mutable; aColor : Color from Draw)
        ---C++: inline
     is static;

  PolesColor (me)  returns Color from Draw
        ---C++: inline
     is static;
    
  Copy(me) returns mutable Drawable3D from Draw
	---Purpose: For variable copy.
  is redefined;
  
      
fields

  drawPoles  : Boolean;
  polesLook  : Color from Draw;

end BezierCurve2d;
