-- File:        SurfacePatch.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSurfacePatch from RWStepGeom

	---Purpose : Read & Write Module for SurfacePatch

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SurfacePatch from StepGeom,
     EntityIterator from Interface

is

	Create returns RWSurfacePatch;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable SurfacePatch from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : SurfacePatch from StepGeom);

	Share(me; ent : SurfacePatch from StepGeom; iter : in out EntityIterator);

end RWSurfacePatch;
