-- File:        VertexLoop.cdl
-- Created:     Mon Dec  4 12:02:33 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWVertexLoop from RWStepShape

	---Purpose : Read & Write Module for VertexLoop

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     VertexLoop from StepShape,
     EntityIterator from Interface

is

	Create returns RWVertexLoop;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable VertexLoop from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : VertexLoop from StepShape);

	Share(me; ent : VertexLoop from StepShape; iter : in out EntityIterator);

end RWVertexLoop;
