-- File:	IGESBasic_ToolGroupWithoutBackP.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolGroupWithoutBackP  from IGESBasic

    ---Purpose : Tool to work on a GroupWithoutBackP. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses GroupWithoutBackP from IGESBasic,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolGroupWithoutBackP;
    ---Purpose : Returns a ToolGroupWithoutBackP, ready to work


    ReadOwnParams (me; ent : mutable GroupWithoutBackP;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : GroupWithoutBackP;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : GroupWithoutBackP;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a GroupWithoutBackP <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable GroupWithoutBackP) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a GroupWithoutBackP
    --           (Null Elements are removed from list)

    DirChecker (me; ent : GroupWithoutBackP) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : GroupWithoutBackP;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : GroupWithoutBackP; entto : mutable GroupWithoutBackP;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : GroupWithoutBackP;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolGroupWithoutBackP;
