-- File:	RWStepFEA_RWFeaModel.cdl
-- Created:	Thu Dec 12 17:51:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFeaModel from RWStepFEA

    ---Purpose: Read & Write tool for FeaModel

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FeaModel from StepFEA

is
    Create returns RWFeaModel from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FeaModel from StepFEA);
	---Purpose: Reads FeaModel

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FeaModel from StepFEA);
	---Purpose: Writes FeaModel

    Share (me; ent : FeaModel from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFeaModel;
