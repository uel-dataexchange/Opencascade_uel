-- File:	Prs2d_DrawSymbol.cdl
-- Created:	October 2000
-- Author:	TCL

---Copyright:	Matra Datavision 2000

class DrawSymbol from Prs2d inherits Line from Graphic2d

	---Purpose: The primitive symbol for drawing

uses

	Drawer		    from Graphic2d,
	GraphicObject	from Graphic2d, 
    TypeOfSymbol    from Prs2d,
    FStream         from Aspect

raises

	SymbolDefinitionError from Prs2d

is
	-------------------------
	-- Category: Constructor
	-------------------------

	Create( aGO       : GraphicObject from Graphic2d;
		    aSymbType : TypeOfSymbol  from Prs2d;
		    aX, aY    : Real          from Standard;
		    aWidth    : Real          from Standard = 10.0;
		    aHeight   : Real          from Standard = 10.0;
		    anAngle   : Real          from Standard = 0.0 )
	 returns mutable DrawSymbol from Prs2d 
     raises SymbolDefinitionError from Prs2d;

	---Level: Public
	---Purpose: Creates the predefined marker index <anIndex> 
	--	    at position <aX>, <aY> and size <aWidth>,<aHeight>.
    ---Category: Constructor
	---Purpose:  Trigger  -   Raises SymbolDefinitionError if the
	--	    symbol type isn't defined,
	--      or the symbol size < aWidth, aHeight > is null.

	----------------------------------------------------
	-- Category: Draw and Pick
	----------------------------------------------------

	Draw( me: mutable; aDrawer: Drawer from Graphic2d ) is static protected;
	---Level: Internal
	---Purpose: Draws the symbol <me>.

	Pick( me : mutable; 
          X, Y       : ShortReal from Standard;
		  aPrecision : ShortReal from Standard;
		  aDrawer    : Drawer from Graphic2d ) returns Boolean from Standard
	  is static protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the symbol <me> is picked,
	--	    Standard_False if not.
	--  Warning: Checks only if the point <X>, <Y> is in the
	--	    boundary rectangle of <me>

   Save( me; aFStream: in out FStream from Aspect ) is virtual;

fields

	myTypeSymb : TypeOfSymbol from Prs2d;
	myX        : ShortReal from Standard;
	myY        : ShortReal from Standard;
	myWidth    : ShortReal from Standard;
	myHeight   : ShortReal from Standard;
	myAngle    : ShortReal from Standard;

end Marker from Graphic2d;
