-- File:	StepRepr_ItemDefinedTransformation.cdl
-- Created:	Wed Mar 26 14:38:45 1997
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


class ItemDefinedTransformation  from StepRepr    inherits TShared

    ---Purpose : Added from StepRepr Rev2 to Rev4

uses
     HAsciiString from TCollection,
     RepresentationItem from StepRepr

is

    Create returns mutable ItemDefinedTransformation;

    Init (me : mutable;
    	  aName : HAsciiString from TCollection;
	  aDescription : HAsciiString from TCollection;
	  aTransformItem1 : RepresentationItem from StepRepr;
	  aTransformItem2 : RepresentationItem from StepRepr);

    SetName (me : mutable; aName : HAsciiString from TCollection);
    Name    (me) returns HAsciiString from TCollection;

    SetDescription (me : mutable; aDescription : HAsciiString from TCollection);
    Description    (me) returns HAsciiString from TCollection;

    SetTransformItem1 (me : mutable; aItem : RepresentationItem from StepRepr);
    TransformItem1    (me) returns RepresentationItem;

    SetTransformItem2 (me : mutable; aItem : RepresentationItem from StepRepr);
    TransformItem2    (me) returns RepresentationItem;

fields

    theName : HAsciiString from TCollection;
    theDescription : HAsciiString from TCollection;
    theTransformItem1 : RepresentationItem from StepRepr;
    theTransformItem2 : RepresentationItem from StepRepr;

end ItemDefinedTransformation;
