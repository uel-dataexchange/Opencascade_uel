-- File:        CsgSelect.cdl
-- Created:     Fri Dec  1 11:11:10 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class CsgSelect from StepShape 

    -- inherits SelectType from StepData

	-- <CsgSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : BooleanResult, CsgPrimitive

uses

	BooleanResult,
	CsgPrimitive
is

	Create returns CsgSelect;
	---Purpose : Returns a CsgSelect SelectType

    	SetTypeOfContent(me : in out; aTypeOfContent : Integer);

	TypeOfContent(me) returns Integer;
	--        1 -> BooleanResult
	--        2 -> CsgPrimitive
	--        0 else
	
	BooleanResult (me) returns any BooleanResult;
	---Purpose : returns Value as a BooleanResult (Null if another type)

    	SetBooleanResult (me : in out;aBooleanResult : BooleanResult from StepShape);
	
	CsgPrimitive (me) returns CsgPrimitive;
	---Purpose : returns Value as a CsgPrimitive (Null if another type)

    	SetCsgPrimitive (me : in out; aCsgPrimitive : CsgPrimitive from StepShape);
	
fields

    theBooleanResult : BooleanResult from StepShape;
    theCsgPrimitive  : CsgPrimitive  from StepShape;  -- a Select Type
    theTypeOfContent : Integer       from Standard;

end CsgSelect;

