-- File:	RWStepShape_RWEdgeBasedWireframeShapeRepresentation.cdl
-- Created:	Fri Dec 28 16:02:01 2001 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWEdgeBasedWireframeShapeRepresentation from RWStepShape

    ---Purpose: Read & Write tool for EdgeBasedWireframeShapeRepresentation

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    EdgeBasedWireframeShapeRepresentation from StepShape

is
    Create returns RWEdgeBasedWireframeShapeRepresentation from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : EdgeBasedWireframeShapeRepresentation from StepShape);
	---Purpose: Reads EdgeBasedWireframeShapeRepresentation

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: EdgeBasedWireframeShapeRepresentation from StepShape);
	---Purpose: Writes EdgeBasedWireframeShapeRepresentation

    Share (me; ent : EdgeBasedWireframeShapeRepresentation from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWEdgeBasedWireframeShapeRepresentation;
