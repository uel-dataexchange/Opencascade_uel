
--Copyright:      Matra Datavision 1992,1993

-- File:          OSD_SharedMemory.cdl
-- Created:       Fri 21 1992
-- Author:        Stephan GARNAUD (ARM)
--                <sga@sparc4>



class SharedMemory from OSD 

   ---Purpose: IPC Tools -Shared Memory
   --          This is a low level interface for communications.
   --          Using shared memory, processes can use a common area to
   --          communicate.
   --          You can create and delete a shared memory.

uses Error, AsciiString from TCollection
raises ConstructionError, NullObject, OSDError, ProgramError
   

is
  Create returns SharedMemory;
    ---Purpose: Allocates room for shared memory name.
    --          This is to be used with 'Open'.
    --          In this case, the process is a client of shared memory.
    ---Level: Advanced

  Create (Name : AsciiString ; size : Integer) returns SharedMemory
    ---Purpose: Instantiates SharedMemory object with parameters.
    --          A name to make sure shared memory is unique and a size in
    --          bytes for the size of shared memory.
    --
    --          Raises ConstructionError when the name contains characters 
    --          not in range of ' '...'~'.
    --          Raises ProgramError when the size given is negative or null.
    --          This is for a server process.
    --          
    ---Level: Advanced
    raises ConstructionError, ProgramError;

  Build (me : in out)  is static;
    ---Purpose: Creates a shared memory in the system
    --          This is for a server process.
    ---Level: Advanced

  Open (me : in out ; Name : AsciiString ; size : Integer)
    ---Purpose: Opens a shared memory
    --          Raises ConstructionError when the name contains characters 
    --          not in range of ' '...'~'.
    --          Raises ProgramError when the size given is negative or null.
    --          This is for a server process.
    --          
    ---Level: Advanced
    raises ConstructionError, ProgramError is static;

  Delete (me : in out)
    ---Purpose: Removes a shared memory access.
    --          This is used only by a server process !
    ---Level: Advanced
    raises ProgramError is static;

  GiveAddress (me) returns Address
    ---Purpose: Returns address of shared memory.
    --          Raises NullObject when the Shared Memory is not created.
    ---Level: Advanced
    raises NullObject is static;

  Failed (me) returns Boolean is static;
    ---Purpose: Returns TRUE if an error occurs
    ---Level: Advanced

  Reset (me : in out) is static;
    ---Purpose: Resets error counter to zero
    ---Level: Advanced
      
  Perror (me : in out)
    ---Purpose: Raises OSD_Error
    ---Level: Advanced
    raises OSDError is static;

 Error (me) returns Integer is static;
   ---Purpose: Returns error number if 'Failed' is TRUE.
    ---Level: Advanced

fields
   myId : Integer;     -- Shared memory ID
   myAddress    : Address;
   myName : AsciiString;   
   mySize : Integer;
   myError : Error;
end SharedMemory from OSD;

