-- File:        DraughtingPreDefinedColour.cdl
-- Created:     Mon Dec  4 12:02:25 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWDraughtingPreDefinedColour from RWStepVisual

	---Purpose : Read & Write Module for DraughtingPreDefinedColour

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     DraughtingPreDefinedColour from StepVisual

is

	Create returns RWDraughtingPreDefinedColour;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable DraughtingPreDefinedColour from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : DraughtingPreDefinedColour from StepVisual);

end RWDraughtingPreDefinedColour;
