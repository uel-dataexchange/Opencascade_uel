
-- File:	Graphic2d_Text.cdl
-- Created:	Tue Jun 22 16:36:51 1993
-- Author:	Jean Louis FRENKEL, Gerard GRAS
--		<jlf@stylox>
-- Modified: TCL G002A, 28-11-00, new inquire methods GetText() and GetType()

---Copyright:	 Matra Datavision 1993

class Text from Graphic2d inherits Primitive from Graphic2d

	---Version:

	---Purpose: The primitive Text

	---Keywords: Primitive, Text
	---Warning:
	---References:

uses
	Drawer		from Graphic2d,
	GraphicObject	from Graphic2d,
	TypeOfAlignment	from Graphic2d,
	PlaneAngle	from Quantity,
	Length		from Quantity,
	Factor		from Quantity,
	ExtendedString	from TCollection,
	TypeOfText	from Aspect,
	FStream		from Aspect,
	IFStream	from Aspect



is
	-------------------------
	-- Category: Constructors
	-------------------------

	Create (aGraphicObject: GraphicObject from Graphic2d;
		aText: ExtendedString from TCollection;
		X, Y: Real from Standard;
		anAngle: PlaneAngle from Quantity = 0.0;
		aType: TypeOfText from Aspect = Aspect_TOT_SOLID;
		aScale: Factor from Quantity = 1.0)
	returns mutable Text from Graphic2d;
	---Level: Public
	---Purpose: Creates a text in a graphic object <aGraphicObject>
	--	    The text is <aText>.
	--	    The reference point is <X>, <Y>.
	--	    The orientation angle is <anAngle>.
	--	    The type of text is <aType> and must be one of :
	--		Aspect_TOT_SOLID,
	--		Aspect_TOT_OUTLINE,
	--	    The scale factor apply to the original font size,
	--	    Angles are measured counterclockwise with 0 radian
	--	    at 3 o'clock.
	--  Warning: a text can be orientable,slantable,zoomable or outlinable
	-- only when this options are enable regardless of the graphic driver.
	-- i.e: Xw driver does not,but Xdps or PS driver does.
	---Category: Constructors

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetFontIndex (me:mutable; anIndex: Integer from Standard = 0)
	is static;
	---Level: Public
	---Purpose: Sets the font index for the text <me>.
        --  Warning: Note that the index 0 can be undefined as a FontMapEntry,
        --        in this case the default system text font is taken.

	SetSlant (me: mutable; aSlant: PlaneAngle from Quantity = 0.0)
	is static;
	---Level: Public
	---Purpose: Sets the slant angle of the text <me>.

        SetZoomable (me: mutable; aFlag: Boolean from Standard = Standard_True)
        is static;
	---Level: Public
        ---Purpose: The text <me> follows the scale factor of the view
        --          if the flag is Standard_True.
        ---Category: Zoom management

	SetOffset (me: mutable; aDx: Real from Standard = 0.0;
				aDy: Real from Standard = 0.0)
        is static;
	---Level: Public
	---Purpose: Sets the Device space offset of the text <me>.

	SetUnderline (me: mutable; 
		isUnderlined: Boolean from Standard = Standard_False)
        is static;
	---Level: Public
	---Purpose: Enable/Disable text underline.

        SetAlignment (me:mutable; anAlignment: TypeOfAlignment from Graphic2d =
                                                        Graphic2d_TOA_LEFT)
        is static;
        ---Level: Public
        ---Purpose: Sets the  text alignment.

	Fit (me:mutable; aWidth,aHeight: Length from Quantity;
			 Adjust: Boolean from Standard = Standard_True; 
			 Expand: Boolean from Standard = Standard_True) 
			returns Boolean from Standard is virtual;
        ---Level: Public
        ---Purpose: Compute text size depending of a required bounding box,
	--	    Adjust the text position depending of the text origine
	--	    and base line if "Adjust" is TRUE,
	--	    Expand the text when the Width is smaller that the
	--	    Fit Width if "Expand" is TRUE.
        --          and returns Standard_True if the current Driver used is 
	--	    enable to fit the text size.
	--  Warning: The fit computation is apply only if the corresponding
	-- dimension is > 0.

	Trunc (me:mutable; aWidth: Length from Quantity)
			returns Boolean from Standard is virtual;
        ---Level: Public
        ---Purpose: Trunc the text when the Width of the text is greater
	--	    that the defined Width Max,
        --          and returns Standard_True if the current Driver used is 
	--	    enable to trunc the text size.

	--------------------------
	-- Category: Draw and Pick
	--------------------------

	Draw (me : mutable; aDrawer: Drawer from Graphic2d)
	is virtual protected;
	---Level: Internal
	---Purpose: Draws the text <me>.

	Pick (me : mutable; X, Y: ShortReal from Standard;
		aPrecision: ShortReal from Standard;
		aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard
	is virtual protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the text <me> is picked,
	--	    Standard_False if not.

        ----------------------------
        -- Category: Inquire methods
        ----------------------------
 
    IsZoomable (me)
                returns Boolean from Standard is static;
    ---Level: Public 
    ---Purpose: Returns Standard_True if the Text <me> follows
    --          the scale factor of the view.
    ---Category: Zoom management

	IsUnderlined (me) returns Boolean from Standard is static;
        ---Level: Public 
        ---Purpose: Returns Standard_True if the Text <me> is underlined.

	TextSize (me; aWidth,aHeight: out Length from Quantity)
                returns Boolean from Standard is static;
        ---Level: Public 
        ---Purpose: Returns Standard_True if the current Driver used is enabled
	--	   to get the right size in the 
	--	   world size parameter <aWidth>,<aHeight> 
	--	   depending of the attributes of the text and the current scale
	--	   of the view.
        ---Category: Text management

	TextSize (me; aWidth,aHeight,anXoffset,anYoffset: out Length from Quantity)
                returns Boolean from Standard is virtual;
        ---Level: Public 
        ---Purpose: Returns Standard_True if the current Driver used is enabled
	--	   to get the right size and text offsets in the 
	--	   world size parameter <aWidth>,<aHeight>,<anXoffset>,<anYoffset> 
	--	   depending of the attributes of the text and the current scale
	--	   of the view.
	--	    NOTE that the text offsets defines the relative position of the 
	--	   of the text string origin from the lower left corner of the text  
	--	   boundary limits.
        ---Category: Text management

	Position (me; X,Y: out Length from Quantity) is static;
        ---Level: Public 
        ---Purpose: Returns the text position.

	Offset (me; X,Y: out Real from Standard) is static;
        ---Level: Public 
        ---Purpose: Returns the text Offset.

	Slant (me) returns PlaneAngle from Quantity is static;
        ---Level: Public 
        ---Purpose: Returns the text slant.

	Angle (me) returns PlaneAngle from Quantity is static;
        ---Level: Public 
        ---Purpose: Returns the text orientation.
                                           
	FontIndex (me) returns Integer from Standard is static;
        ---Level: Public 
        ---Purpose: Returns the text font index.

	Scale (me) returns Factor from Quantity is static;
        ---Level: Public 
        ---Purpose: Returns the text scale.

    Alignment (me) returns TypeOfAlignment from Graphic2d is static;
        ---Level: Public
        ---Purpose: Returns the text alignment.

    GetText( me ) returns ExtendedString from TCollection;
    ---Level: Public
    ---Purpose: Returns the text string

    GetType( me ) returns TypeOfText from Aspect;
    ---Level: Public
    ---Purpose: Returns the type text

    ----------------------------
    -- Category: Private methods
    ----------------------------

	ComputeMinMax (me : mutable) 
		returns Boolean from Standard is redefined virtual protected;
        ---Level: Internal
        ---Purpose: Computes the MinMax of the text if possible.

	----------------------------------------------------------------------

	Save( me; aFStream: in out FStream from Aspect ) is virtual;
--	Retrieve( me; aIFStream: in out IFStream from AIS2D ) is virtual;

fields

	myFontIndex:    Integer from Standard is protected;

	myX,myDx:	    ShortReal from Standard is protected;
	myY,myDy:	    ShortReal from Standard is protected;
	myAngle:	    ShortReal from Standard is protected;
	myType:		    TypeOfText from Aspect is protected;
	myText:		    ExtendedString from TCollection is protected;
	myAdjustFlag:   Boolean from Standard is protected;

	myDeltax:	    ShortReal from Standard is protected;
	myDeltay:	    ShortReal from Standard is protected;
	mySlant:	    ShortReal from Standard is protected;
	myIsZoomable:   Boolean from Standard is protected;
	myIsUnderlined:	Boolean from Standard is protected;
	myHScale:	    Factor from Quantity is protected;
	myWScale:	    Factor from Quantity is protected;
	myAlignment:	TypeOfAlignment from Graphic2d is protected;

end Text from Graphic2d;
