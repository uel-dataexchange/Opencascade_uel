-- File:        TextLiteral.cdl
-- Created:     Mon Dec  4 12:02:32 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWTextLiteral from RWStepVisual

	---Purpose : Read & Write Module for TextLiteral

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     TextLiteral from StepVisual,
     EntityIterator from Interface

is

	Create returns RWTextLiteral;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable TextLiteral from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : TextLiteral from StepVisual);

	Share(me; ent : TextLiteral from StepVisual; iter : in out EntityIterator);

end RWTextLiteral;
