-- File:	RWStepFEA_RWFreedomsList.cdl
-- Created:	Sat Dec 14 11:02:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFreedomsList from RWStepFEA

    ---Purpose: Read & Write tool for FreedomsList

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FreedomsList from StepFEA

is
    Create returns RWFreedomsList from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FreedomsList from StepFEA);
	---Purpose: Reads FreedomsList

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FreedomsList from StepFEA);
	---Purpose: Writes FreedomsList

    Share (me; ent : FreedomsList from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFreedomsList;
