-- File:	BOP_WireEdgeSet.cdl
-- Created:	Wed Jun 16 11:52:45 1993
-- Author:	Jean Yves LEBEY
--		<jyl@zerox>
---Copyright:	 Matra Datavision 1993

class WireEdgeSet from BOP inherits ShapeSet from BOP

    ---Purpose: The class containing data and methods  
    --          for a set of edges and wires
    --
    -- Bound is a wire,  
    -- Boundelement is an edge.
    --
    -- The ShapeSet stores :
    --  - a list of wire (bounds),
    --  - a list of edge (boundelements) to start reconstructions,
    --  - a map of vertex giving the list of edge incident to a vertex.

uses

    Orientation from TopAbs, 
    
    Shape  from TopoDS,
    Face   from TopoDS,
    Edge   from TopoDS,
    Vertex from TopoDS,
    
    ListOfShape from TopTools, 
    
    Pnt2d from gp,
    Vec2d from gp
   
    
is
    Create   
    	returns WireEdgeSet from BOP; 
    	---Purpose:  
    	--- Empty constructor; 
    	---
    Create  (F:  Face from TopoDS) 
    	returns WireEdgeSet from BOP;
    	---Purpose:  
    	--- Creates a WES to build edges connected by vertices
    	--- on face F. Edges of the WireEdgeSet must have a representation
    	--- on surface of face F.
    	---
    Initialize(me:out; 
    	    F:  Face from TopoDS);   
    	---Purpose:  
    	--- Initialize a WES to build edges connected by vertices
    	--- on face F. Edges of the WireEdgeSet must have a representation
    	--- on surface of face F. 
    	---
    Face(me)  
    	returns Face from TopoDS;
    	---C++: return const & 
    	---Purpose:   
    	--- Selector 
    	---
    AddShape(me:out; 
    	    S:Shape from TopoDS)  
    	is redefined;
    	---Purpose:    
    	--- See  in  base  class,  please  
    	---
    AddStartElement(me:out; 
    	    S:Shape from TopoDS)  
    	is redefined;
    	---Purpose:    
    	--- See  in  base  class,  please  
    	---
    AddElement(me:out; 
    	    S:Shape from TopoDS)  
    	is redefined;
    	---Purpose:    
    	--- See  in  base  class,  please  
    	---
    InitNeighbours(me:out; 
    	    E:Shape from TopoDS)  
    	is redefined; 
    	---Purpose:  
    	--- Internal  usage 
    	---
    FindNeighbours(me:out)  
    	is redefined;
    	---Purpose:
    	--- Build the list of neighbour edges of edge myCurrentShape
    	--- Initialize iterator of neighbour edges to edge myCurrentShape
    	---
    MakeNeighboursList(me:out; 
    	    	       E,V:Shape from TopoDS)  
    	returns ListOfShape from TopTools  
    	is redefined;
    	---C++: return const &
   
    VertexConnectsEdges(me; 
    	    V,E1,E2:Shape from TopoDS; 
    	    O1,O2:out Orientation from TopAbs)
    	returns Boolean from Standard 
    	is private;
    	---Purpose: 
    	--- Indicates whether vertex V is a good connexity vertex between
    	--- edges E1 and E2.
    	--- i.e, returns True if V is shared by E1 and E2 and if V has different 
    	--- orientations on E1 and E2.
    	--- If V is shared by E1 and E2, returns the orientation of V on E1 and E2
	---

    VertexConnectsEdgesClosing(me; 
    	    V,E1,E2:Shape from TopoDS)  
    	returns Boolean from Standard 
    	is private;
    	---Purpose:  
    	--- Internal  usage 
    	---
    NbClosingShapes(me; 
    	    L:ListOfShape from TopTools)  
    	returns Integer from Standard  
    	is private;
    	---Purpose:  
    	--- Internal  usage 
    	---
    LocalD1(me; 
    	    F :  Face from  TopoDS; 
    	    E :  Edge from  TopoDS;  
    	    V :  Vertex from TopoDS; 
    	    P2:  out Pnt2d from gp; 
    	    V2:  out Vec2d from gp)  
    	is private;
    	---Purpose:  
    	--- Internal  usage 
    	---
    IsClosed(me; 
    	    E:Shape from TopoDS) 
    	 returns Boolean from Standard 
    	 is private;
    	---Purpose:  
    	--- indicates if the edge <E> is a closing edge of myFace
    	--- Internal  usage 
    	---
    IsUClosed(me; 
    	    E:Shape from TopoDS)  
    	returns Boolean from Standard  
    	is private;
    	---Purpose:  
    	--- indicates if the edge <E> is a closing edge on U of myFace
    	--- Internal  usage 
    	---
    IsVClosed(me; 
    	    E:Shape from TopoDS)  
    	returns Boolean from Standard  
    	is private;
    	---Purpose:  
    	--- indicates if the edge <E> is a closing edge on V of myFace
    	--- Internal  usage 
    	---
    IsUVISO(myclass; 
    	    E:Edge from TopoDS; 
    	    F:Face from TopoDS; 
    	    uiso,viso:out Boolean from Standard);
    	---Purpose:  
    	--- Internal  usage 
    	---

    RemoveEdgeFromWES  (me:out; 
    	    aE : Edge from TopoDS);
    	---Purpose:  
    	--- Removes the edge aE from the WES      
    	---
    KeptTwice(me; 
    	    aE : Edge from  TopoDS) 
    	returns Boolean from Standard;   
    	---Purpose:  
    	--- Returns TRUE if the edge aE has been kept twice 
    	--- in  the WES      
    	---
    
fields

    myFace:Face from TopoDS;
    myDEBVertexIndex:Integer from Standard;
    
end WireEdgeSet from BOP;
