-- File:        GeometricSetSelect.cdl
-- Created:     Fri Dec  1 11:11:11 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class GeometricSetSelect from StepShape inherits SelectType from StepData

	-- <GeometricSetSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : Point, Curve, Surface

uses

	Point   from StepGeom,
	Curve   from StepGeom,
	Surface from StepGeom
is

	Create returns GeometricSetSelect;
	---Purpose : Returns a GeometricSetSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a GeometricSetSelect Kind Entity that is :
	--        1 -> Point
	--        2 -> Curve
	--        3 -> Surface
	--        0 else

	Point (me) returns any Point;
	---Purpose : returns Value as a Point (Null if another type)

	Curve (me) returns any Curve;
	---Purpose : returns Value as a Curve (Null if another type)

	Surface (me) returns any Surface;
	---Purpose : returns Value as a Surface (Null if another type)


end GeometricSetSelect;

