-- File:	MakeMirror.cdl
-- Created:	Tue Sep  1 15:33:36 1992
-- Author:	Remi GILET
--		<reg@sdsun1>
---Copyright:	 Matra Datavision 1992

class MakeMirror

from gce

    ---Purpose: This class mplements elementary construction algorithms for a
    -- symmetrical transformation in 3D space about a point,
    -- axis or plane. The result is a gp_Trsf transformation.
    -- A MakeMirror object provides a framework for:
    -- -   defining the construction of the transformation,
    -- -   implementing the construction algorithm, and
    -- -   consulting the result.
 

uses Pnt  from gp,
     Ax1  from gp,
     Ax2  from gp,
     Dir  from gp,
     Pln  from gp,
     Lin  from gp,
     Trsf from gp,
     Real from Standard
     
is

Create(Point : Pnt from gp) returns MakeMirror;
    ---Puprose: Makes a symmetry transformation of center <Point>.

Create(Axis : Ax1 from gp) returns MakeMirror;
    ---Puprose: Makes a symmetry transformation of axis <Axis>.

Create(Line : Lin from gp) returns MakeMirror;
    ---Puprose: Makes a symmetry transformation of axis <Line>.

Create(Point : Pnt from gp;
       Direc : Dir from gp) returns MakeMirror;
    ---Purpose: Makes a symmetry transformation af axis defined by 
    --          <Point> and <Direc>.

Create(Plane : Pln from gp) returns MakeMirror;
    ---Purpose: Makes a symmetry transformation of plane <Plane>.

Create(Plane : Ax2 from gp) returns MakeMirror;
    ---Purpose: Makes a symmetry transformation of plane <Plane>.

Value(me) returns Trsf from gp
    is static;
    ---C++: return const&
    ---Purpose: Returns the constructed transformation.
    
Operator(me) returns Trsf from gp
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator gp_Trsf() const;"

fields

    TheMirror : Trsf from gp;

end MakeMirror;

