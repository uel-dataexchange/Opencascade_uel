-- File:	BRepSweep_Trsf.cdl
-- Created:	Tue Jun  8 15:43:21 1993
-- Author:	Laurent BOURESCHE
--		<lbo@phobox>
---Copyright:	 Matra Datavision 1993


deferred class Trsf from BRepSweep inherits NumLinearRegularSweep 
    	    	    	    	    	    from BRepSweep

	---Purpose: This class is inherited from NumLinearRegularSweep
	--          to  implement the  simple   swept primitives built
	--          moving a Shape with a Trsf.  It  often is possible
	--          to  build  the constructed subshapes  by  a simple
	--          move of the  generating subshapes (shared topology
	--          and geometry).   So two  ways of construction  are
	--          proposed : 
	--          
    	--
	--          - sharing  basis elements  (the generatrice can be
	--          modified , for  exemples  PCurves can be added  on
	--          faces);
    	--
	--          - copying everything.


uses

    Builder from BRep,
    Shape from TopoDS,
    NumShape from Sweep,
    Location from TopLoc,
    Orientation from TopAbs
    
is

    Delete(me:out) is redefined;
    ---C++: alias "Standard_EXPORT virtual ~BRepSweep_Trsf(){Delete() ; }"
    
    Initialize(aBuilder  : Builder from BRep;
               aGenShape : Shape from TopoDS;
    	       aDirWire  : NumShape from Sweep;
    	       aLocation : Location from TopLoc;
    	       aCopy     : Boolean from Standard);
	---Purpose: Initialize  the Trsf BrepSweep, if  aCopy  is true
	--          the  basis elements  are    shared  as   often  as
	--          possible, else everything is copied.
    	--          

    Init(me : in out)
    	---Purpose: ends  the  construction  of the   swept  primitive
    	--          calling the virtual geometric functions that can't
    	--          be called in the initialize.
    is static;

    Process (me    : in out;
    	     aGenS : Shape from TopoDS;
    	     aDirV : NumShape from Sweep) 
    returns Boolean from Standard
    	---Purpose: function called to analize the way of construction
    	--          of the shapes generated by aGenS and aDirV.
    is static;

    -- """"""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""
    --  Deferred Methods supporting the creation of the geometric part.
    -- """"""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""
    
    MakeEmptyVertex(me    : in out; 
    	    	    aGenV : Shape from TopoDS; 
    	    	    aDirV : NumShape from Sweep)
    returns Shape from TopoDS 
	---Purpose: Builds the vertex addressed by [aGenV,aDirV], with its
	--          geometric part, but without subcomponents.
    is deferred;
    
    MakeEmptyDirectingEdge(me    : in out; 
    	    	    	   aGenV : Shape from TopoDS; 
    	    	    	   aDirE : NumShape from Sweep)
    returns Shape from TopoDS
	---Purpose: Builds the edge addressed by [aGenV,aDirE], with its
	--          geometric part, but without subcomponents.
    is deferred;
    
    MakeEmptyGeneratingEdge(me    : in out; 
    	    	    	    aGenE : Shape from TopoDS; 
    	    	    	    aDirV : NumShape from Sweep)
    returns Shape from TopoDS
	---Purpose: Builds the edge addressed by [aGenE,aDirV], with its
	--          geometric part, but without subcomponents.
    is deferred;
    
    SetParameters(me         : in out; 
    	    	  aNewFace   : Shape from TopoDS; 
    	      	  aNewVertex : in out Shape from TopoDS;
    	    	  aGenF      : Shape from TopoDS; 
    	    	  aGenV      : Shape from TopoDS;
    	    	  aDirV      : NumShape from Sweep)
	---Purpose: Sets the  parameters of the new  vertex  on the new
	--          face. The new face and  new vertex where generated
	--          from aGenF, aGenV and aDirV .
    is deferred;
    
    SetDirectingParameter(me         : in out; 
    	    	          aNewEdge   : Shape from TopoDS; 
    	    	    	  aNewVertex : in out Shape from TopoDS;
    	    	          aGenV      : Shape from TopoDS;
    	    	          aDirE      : NumShape from Sweep; 
    	    	    	  aDirV      : NumShape from Sweep)
	---Purpose: Sets the  parameter of the new  vertex  on the new
	--          edge. The new edge and  new vertex where generated
	--          from aGenV aDirE, and aDirV.
    is deferred;

    SetGeneratingParameter(me         : in out; 
    	    	    	   aNewEdge   : Shape from TopoDS; 
                           aNewVertex : in out Shape from TopoDS;
    	    	    	   aGenE      : Shape from TopoDS; 
                           aGenV      : Shape from TopoDS;
    	    	    	   aDirV      : NumShape from Sweep)
	---Purpose: Sets the  parameter of the new  vertex  on the new
	--          edge. The new edge and  new vertex where generated
	--          from aGenE, aGenV and aDirV .
    is deferred;

    MakeEmptyFace(me       : in out; 
    	    	  aGenS    : Shape from TopoDS; 
    	    	  aDirS    : NumShape from Sweep)
    returns Shape from TopoDS
	---Purpose: Builds  the face addressed  by [aGenS,aDirS], with
	--          its geometric part, but without subcomponents. The
	--          couple aGenS, aDirS can be  a "generating face and
	--          a  directing vertex" or "a   generating edge and a
	--          directing  edge".
    is deferred;
    
    SetPCurve(me       : in out;
 	      aNewFace : Shape from TopoDS; 
              aNewEdge : in out Shape from TopoDS;
	      aGenF    : Shape from TopoDS; 
              aGenE    : Shape from TopoDS;
	      aDirV    : NumShape from Sweep;
              orien    : Orientation from TopAbs)
	 ---Purpose: Sets the PCurve for a new edge on a new face. The
	 --          new edge and  the  new face were generated  using
	 --          aGenF, aGenE and aDirV.
    is deferred;
    
    SetGeneratingPCurve(me       : in out;
    	    	    	aNewFace : Shape from TopoDS; 
                        aNewEdge : in out Shape from TopoDS;
			aGenE    : Shape from TopoDS; 
                        aDirE    : NumShape from Sweep;
			aDirV    : NumShape from Sweep;
                        orien    : Orientation from TopAbs)

	 ---Purpose: Sets the PCurve for a new edge on a new face. The
	 --          new edge and  the  new face were generated  using
	 --          aGenE, aDirE and aDirV.
    is deferred;
    	    
    SetDirectingPCurve(me       : in out;
    	    	       aNewFace : Shape from TopoDS; 
                       aNewEdge : in out Shape from TopoDS;
		       aGenE    : Shape from TopoDS; 
		       aGenV    : Shape from TopoDS; 
                       aDirE    : NumShape from Sweep;
                       orien    : Orientation from TopAbs)

	 ---Purpose: Sets the PCurve for a new edge on a new face. The
	 --          new edge and  the  new face were generated  using
	 --          aGenE, aDirE and aGenV.
    is deferred;
    
    GGDShapeIsToAdd (me;
    	    	     aNewShape    : Shape from TopoDS;
    	    	     aNewSubShape : Shape from TopoDS;
      	    	     aGenS        : Shape from TopoDS;
		     aSubGenS     : Shape from TopoDS;
    	    	     aDirS        : NumShape from Sweep)
    returns Boolean from Standard
	---Purpose: Returns   true   if  aNewSubShape    (addressed by
	--          aSubGenS  and aDirS)  must  be added  in aNewShape
	--          (addressed by aGenS and aDirS).
    is deferred;
    
    GDDShapeIsToAdd (me;
    	    	     aNewShape    : Shape from TopoDS;
    	    	     aNewSubShape : Shape from TopoDS;
      	    	     aGenS        : Shape from TopoDS;
    	    	     aDirS        : NumShape from Sweep;
   	    	     aSubDirS     : NumShape from Sweep)
    returns Boolean from Standard
	---Purpose: Returns   true   if  aNewSubShape    (addressed by
	--          aGenS  and aSubDirS)  must  be added  in aNewShape
	--          (addressed by aGenS and aDirS).
    is deferred;

    SeparatedWires  (me;
    	    	     aNewShape    : Shape from TopoDS;
    	    	     aNewSubShape : Shape from TopoDS;
      	    	     aGenS        : Shape from TopoDS;
		     aSubGenS     : Shape from TopoDS;
    	    	     aDirS        : NumShape from Sweep)
    returns Boolean from Standard
	---Purpose: In  some  particular  cases  the   topology  of  a
	--          generated  face must be  composed  of  independant
	--          closed wires,  in this case  this function returns
	--          true.
    is deferred;
    
    HasShape(me; aGenS : Shape from TopoDS; aDirS : NumShape from Sweep) 
    returns Boolean from Standard
	---Purpose: Returns true   if aDirS   and aGenS  addresses   a
	--          resulting Shape. In some  specific cases the shape
	--          can  be    geometrically   inexsistant,  then this
	--          function returns false.
    is deferred;

    IsInvariant (me; aGenS : Shape from TopoDS)
    returns Boolean from Standard
    	---Purpose: Returns  true if  the geometry   of  aGenS is  not
    	--          modified by the trsf of the BRepSweep Trsf.
    is deferred;


    -- """"""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""
    --  Method coding the continuities on the edges between 2 faces
    -- """"""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""
    SetContinuity(me : in out; 
    	    	  aGenS : Shape from TopoDS; 
    	    	  aDirS : NumShape from Sweep);
       ---Purpose: Called to propagate the continuity of  every vertex
       --          between two edges of the  generating wire  aGenS on
       --          the generated edge and faces.

fields

    myLocation : Location from TopLoc is protected;
    myCopy     : Boolean from Standard is protected;
    
end Trsf from BRepSweep;
