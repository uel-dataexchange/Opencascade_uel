-- File:	MDataStd_IntPackedMapRetrievalDriver_1.cdl
-- Created:	Fri Mar 28 11:31:18 2008
-- Author:	Sergey ZARITCHNY
--		<sergey.zaritchny@opencascade.com>
---Copyright:	Open CasCade SA 2008 


class IntPackedMapRetrievalDriver_1 from MDataStd inherits ARDriver from MDF

	---Purpose: Retrieval  driver of IntPackedMap attribute supporting 
	--          delta mechanism by default

uses
    RRelocationTable from MDF,
    Attribute        from PDF,
    Attribute        from TDF, 
    MessageDriver    from CDM 

is
    Create(theMessageDriver : MessageDriver from CDM)
    returns mutable IntPackedMapRetrievalDriver_1 from MDataStd;
    

    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 1.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type: IntPackedMap_1 from PDataStd.

    NewEmpty (me)  returns mutable Attribute from TDF;


    Paste(me;
    	  Source     :         Attribute from PDF;
    	  Target     : mutable Attribute from TDF;
    	  RelocTable : RRelocationTable  from MDF);



end IntPackedMapRetrievalDriver_1;
