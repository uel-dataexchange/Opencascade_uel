-- File:	BRepLib_FuseEdges.cdl
-- Created:	Mon Sep 10 10:36:48 2007
-- Author:	Igor FEOKTISTOV
--		<ifv@philipox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2007


class FuseEdges from BRepLib 

	---Purpose: This class can detect  vertices in a face that can
	--          be considered useless and then perform the fuse of
	--          the  edges and remove  the  useless vertices.  By
	--          useles vertices,  we mean :
	--            * vertices that  have  exactly two connex edges 
	--            * the edges connex to the vertex must have 
	--              exactly the same 2 connex faces .
	--            * The edges connex to the vertex must have the
	--               same geometric support.

uses
  Shape from TopoDS,
  Vertex from TopoDS,
  Edge from TopoDS,
  ShapeEnum from TopAbs,
  MapOfShape from TopTools,
  ListOfShape from TopTools,
  DataMapOfIntegerListOfShape from TopTools,
  DataMapOfIntegerShape from TopTools,
  DataMapOfShapeShape from TopTools,
  IndexedDataMapOfShapeListOfShape from TopTools,
  IndexedMapOfShape from TopTools

raises
      	ConstructionError from Standard,
        NullObject        from Standard

is
    Create (theShape : Shape from TopoDS;
            PerformNow : Boolean from Standard = Standard_False)
    returns FuseEdges from BRepLib
    raises NullObject        from Standard;
    	---Purpose: Initialise members  and build  construction of map
    	--          of ancestors.

    AvoidEdges (me : in out; theMapEdg : IndexedMapOfShape from TopTools);
        ---Purpose: set edges to avoid being fused 
	 
    --  Modified  by  IFV  19.04.07   
    SetConcatBSpl(me : in out; theConcatBSpl : Boolean from Standard = Standard_True);
        ---Purpose: set mode to enable concatenation G1 BSpline edges in one 
    --  End  Modified  by  IFV  19.04.07   

    Edges (me : in out ; theMapLstEdg : in out DataMapOfIntegerListOfShape from TopTools);
    	---Purpose: returns  all the list of edges to be fused
    	--          each list of the map represent a set of connex edges
    	--          that can be fused.

    ResultEdges (me : in out ; theMapEdg : in out DataMapOfIntegerShape from TopTools);
    	---Purpose: returns all the fused edges. each integer entry in
    	--           the   map  corresponds  to  the  integer   in the
    	--           DataMapOfIntegerListOfShape  we    get in  method
    	--          Edges.   That is to say, to  the list  of edges in
    	--          theMapLstEdg(i) corresponds the resulting edge theMapEdge(i)
    	--          


    Faces (me: in out; theMapFac : in out DataMapOfShapeShape from TopTools); 
    	---Purpose: returns the map of modified faces.

    Shape (me : in out)
    returns Shape from TopoDS
    raises NullObject        from Standard;
    	---Purpose: returns myShape modified with the list of internal
    	--          edges removed from it.
        ---C++: return &

    NbVertices (me : in out)
    returns Integer from Standard
    raises NullObject        from Standard;
    	---Purpose: returns the number of vertices candidate to be removed
    	---C++: return const

    Perform (me : in out);
    ---Purpose: Using  map of list of connex  edges, fuse each list to
    --           one edge and then update myShape


    BuildAncestors (me; S: Shape from TopoDS; TS: ShapeEnum from TopAbs; 
		    TA: ShapeEnum from TopAbs; M: in out IndexedDataMapOfShapeListOfShape from TopTools)
    ---Purpose: build a map of shapes and ancestors, like 
    --          TopExp.MapShapesAndAncestors, but we remove duplicate 
    --          shapes in list of shapes.
    is private;
    
    BuildListEdges (me : in out)
        ---Purpose: Build the all the lists of edges that are to be fused
    is private;
    
    BuildListResultEdges (me : in out)
        ---Purpose: Build result   fused edges according  to  the list
        --          builtin BuildLisEdges
    is private;
    
    BuildListConnexEdge (me : in out; theEdge : Shape from TopoDS; theMapUniq : in out MapOfShape from TopTools;
    	    	    	 theLstEdg : in out ListOfShape from TopTools)
    is private;
    
    NextConnexEdge (me; theVertex : Vertex from TopoDS; theEdge : Shape from TopoDS; 
    	    	    theEdgeConnex : in out Shape from TopoDS)
    returns Boolean from Standard
    is private;
    
    SameSupport (me; E1 : Edge from TopoDS; E2 :Edge from TopoDS)
    returns Boolean from Standard
    is private;
    
    UpdatePCurve (me; theOldEdge : Edge from TopoDS; 
    	    	      theNewEdge : in out Edge from TopoDS; 
		      theLstEdg  : ListOfShape from TopTools)
    returns Boolean from Standard
    is private;
    
    
fields
    myShape           : Shape from TopoDS;
    myShapeDone       : Boolean from Standard;
    myEdgesDone       : Boolean from Standard;
    myResultEdgesDone : Boolean from Standard;
    myMapVerLstEdg    : IndexedDataMapOfShapeListOfShape from TopTools;
    myMapEdgLstFac    : IndexedDataMapOfShapeListOfShape from TopTools;
    myMapLstEdg       : DataMapOfIntegerListOfShape from TopTools;
    myMapEdg          : DataMapOfIntegerShape from TopTools;
    myMapFaces        : DataMapOfShapeShape from TopTools;
    myNbConnexEdge    : Integer from Standard;
    myAvoidEdg        : IndexedMapOfShape from TopTools; 
    --  Modified  by  IFV  19.04.07   
    myConcatBSpl      : Boolean  from  Standard;  --  to enable  concatenation of G1 BSpline 
                                                  --  edges
    
end FuseEdges;
