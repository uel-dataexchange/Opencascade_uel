-- File:	Dynamic_IntegerParameter.cdl
-- Created:	Wed Feb  3 15:49:43 1993
-- Author:	Gilles DEBARBOUILLE
--		<gde@bravox>
---Copyright:	 Matra Datavision 1993



class IntegerParameter from Dynamic

inherits

    Parameter from Dynamic     
    
	---Purpose: This class describes a parameter with an integer 
	--          as its value.

uses
    CString from Standard,
    Integer from Standard,
    OStream from Standard 

is

    Create(aparameter : CString from Standard)
    
    ---Level: Public 
    
    ---Purpose: Creates   an  IntegerParameter  with  <aparameter>  as
    --          identifier.

    returns mutable IntegerParameter from Dynamic;

    Create(aparameter : CString from Standard ; avalue : Integer from Standard) 

    ---Level: Public 
    
    ---Purpose: Creates   an  IntegerParameter  with  <aparameter>  as
    --          identifier and <avalue> as initial value.

    returns mutable IntegerParameter from Dynamic;
    
    Value(me) returns Integer from Standard
    
    ---Level: Public 
    
    ---Purpose: Returns the integer value <thevalue>.
    
    is static;
    
    Value (me : mutable ; avalue : Integer from Standard)
    
    ---Level: Public 
    
    --- Purpose: Sets the field <thevalue> with the integer value <avalue>

    is static;
    
    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Public 
    
    ---Purpose: Useful for debugging.
    
    is redefined;
    
fields

    thevalue : Integer from Standard;

end IntegerParameter;
