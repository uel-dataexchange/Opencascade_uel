-- File:        Invisibility.cdl
-- Created:     Fri Dec  1 11:11:21 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class Invisibility from StepVisual 

inherits TShared from MMgt

uses

	HArray1OfInvisibleItem from StepVisual, 
	InvisibleItem from StepVisual
is

	Create returns mutable Invisibility;
	---Purpose: Returns a Invisibility

	Init (me : mutable;
	      aInvisibleItems : mutable HArray1OfInvisibleItem from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetInvisibleItems(me : mutable; aInvisibleItems : mutable HArray1OfInvisibleItem);
	InvisibleItems (me) returns mutable HArray1OfInvisibleItem;
	InvisibleItemsValue (me; num : Integer) returns InvisibleItem;
	NbInvisibleItems (me) returns Integer;

fields

	invisibleItems : HArray1OfInvisibleItem from StepVisual; -- a SelectType

end Invisibility;
