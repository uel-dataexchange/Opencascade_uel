-- File:	StepRepr_ProductDefinitionShape.cdl
-- Created:	Mon Jul  3 16:29:03 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class ProductDefinitionShape from StepRepr
inherits PropertyDefinition from StepRepr

    ---Purpose: Representation of STEP entity ProductDefinitionShape

uses
    HAsciiString from TCollection,
    CharacterizedDefinition from StepRepr

is
    Create returns ProductDefinitionShape from StepRepr;
	---Purpose: Empty constructor

end ProductDefinitionShape;
