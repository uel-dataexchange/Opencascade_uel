-- File:	RWStepAP214_RWRepItemGroup.cdl
-- Created:	Wed May 10 15:09:08 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWRepItemGroup from RWStepAP214

    ---Purpose: Read & Write tool for RepItemGroup

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    RepItemGroup from StepAP214

is
    Create returns RWRepItemGroup from RWStepAP214;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : RepItemGroup from StepAP214);
	---Purpose: Reads RepItemGroup

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: RepItemGroup from StepAP214);
	---Purpose: Writes RepItemGroup

    Share (me; ent : RepItemGroup from StepAP214;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWRepItemGroup;
