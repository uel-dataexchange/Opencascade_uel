-- File:        BezierSurfaceAndRationalBSplineSurface.cdl
-- Created:     Mon Dec  4 12:02:34 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWBezierSurfaceAndRationalBSplineSurface from RWStepGeom

	---Purpose : Read & Write Module for BezierSurfaceAndRationalBSplineSurface

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     BezierSurfaceAndRationalBSplineSurface from StepGeom,
     EntityIterator from Interface

is

	Create returns RWBezierSurfaceAndRationalBSplineSurface;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable BezierSurfaceAndRationalBSplineSurface from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : BezierSurfaceAndRationalBSplineSurface from StepGeom);

	Share(me; ent : BezierSurfaceAndRationalBSplineSurface from StepGeom; iter : in out EntityIterator);

end RWBezierSurfaceAndRationalBSplineSurface;
