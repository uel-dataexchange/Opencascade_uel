-- File:        IntPatch_HCurve2dTool.cdl
-- Created:	Mon Jul 17 16:25:23 1995
-- Author:	Laurent BUCHARD
---Copyright:	OPEN CASCADE 1995


class HCurve2dTool from IntPatch

uses 
     HCurve2d        from Adaptor2d,
     Array1OfReal    from TColStd,
     Shape           from GeomAbs,
     CurveType       from GeomAbs,
     Vec2d             from gp,
     Pnt2d             from gp,
     Circ2d            from gp,
     Elips2d           from gp,
     Hypr2d            from gp,
     Parab2d           from gp,
     Lin2d             from gp,
     BezierCurve     from Geom2d,
     BSplineCurve    from Geom2d
     
raises
    
    OutOfRange          from Standard,
    NoSuchObject        from Standard,
    DomainError         from Standard
 
is

    --
    --     Global methods - Apply to the whole curve.
    --     
    
    FirstParameter(myclass; C: HCurve2d from Adaptor2d) returns Real
    	---C++: inline
    ;
    

    LastParameter(myclass; C: HCurve2d from Adaptor2d) returns Real
    	---C++: inline    
    ;

    --
    -- Services to break the curves to the expected continuity
    -- 
    --  If  for example you  need the  curve to  be C2  and the method
    --  Continuity   returns you something lower than   C2 (say C1 for
    --  example).
    --  
    --  First  compute the   number  of intervals  with  the requested
    --  continuity with the method  NbIntervals().   Note that if  the
    --  continuity  is higher than the one   you need NbIntervals will
    --  return 1.
    --  
    --  Then you get the parameters  bounding  the intervals with  the
    --  method  Intervals,   using   an array    of  length  at  least
    --  NbIntervals()+1.
    -- 
    -- If you need  to create a curve  with a restricted span you  can
    -- use the method Trim().

    
    Continuity(myclass; C: HCurve2d from Adaptor2d) returns Shape from GeomAbs
	---Purpose: 
	---C++: inline
    ;
    
    NbIntervals(myclass; C: HCurve2d from Adaptor2d; S : Shape from GeomAbs) returns Integer
	---Purpose: Returns  the number  of  intervals for  continuity
	--          <S>. May be one if Continuity(myclass) >= <S>
	---C++: inline
    ;
    
    Intervals(myclass; C: HCurve2d from Adaptor2d; T : in out Array1OfReal from TColStd; 
    	          S : Shape from GeomAbs)
	---Purpose: Stores in <T> the  parameters bounding the intervals
	--          of continuity <S>.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
    raises
    	OutOfRange from Standard
    ---C++: inline
    ;
    
    IsClosed(myclass; C: HCurve2d from Adaptor2d) returns Boolean
    ---C++: inline    
    ;
     
    IsPeriodic(myclass; C: HCurve2d from Adaptor2d) returns Boolean
    ---C++: inline
    ;
    
    Period(myclass; C: HCurve2d from Adaptor2d) returns Real
    raises
    	DomainError from Standard -- if the curve is not periodic
    ---C++: inline	
    ;
     
    Value(myclass; C: HCurve2d from Adaptor2d; U : Real) returns Pnt2d from gp
         --- Purpose : Computes the point of parameter U on the curve.
    ---C++: inline
    ;
    
    D0 (myclass; C: HCurve2d from Adaptor2d; U : Real; P : out Pnt2d from gp)
         --- Purpose : Computes the point of parameter U on the curve.
    ---C++: inline
    ;
    
    D1 (myclass; C: HCurve2d from Adaptor2d; U : Real; P : out Pnt2d from gp ; V : out Vec2d from gp)
         --- Purpose : Computes the point of parameter U on the curve with its
         --  first derivative.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C1.
    ---C++: inline
    ;
    
    D2 (myclass; C: HCurve2d from Adaptor2d; U : Real; P : out Pnt2d from gp; V1, V2 : out Vec2d from gp)
        --- Purpose :
        --  Returns the point P of parameter U, the first and second
        --  derivatives V1 and V2.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C2.
    ---C++: inline
     ;

    D3 (myclass; C: HCurve2d from Adaptor2d; U : Real; P : out Pnt2d from gp; V1, V2, V3 : out Vec2d from gp)
        --- Purpose :
        --  Returns the point P of parameter U, the first, the second 
        --  and the third derivative.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C3.
    ---C++: inline
     ;
        
    DN (myclass; C: HCurve2d from Adaptor2d; U : Real; N : Integer)   returns Vec2d from gp
        --- Purpose :
        --  The returned vector gives the value of the derivative for the 
        --  order of derivation N.
     raises  
    	DomainError from Standard,
        --- Purpose : Raised if the continuity of the current interval
        --  is not CN.
        OutOfRange from Standard
        --- Purpose : Raised if N < 1.            
    ---C++: inline
     ;

    Resolution(myclass; C: HCurve2d from Adaptor2d; R3d : Real) returns Real
         ---Purpose :  Returns the parametric  resolution corresponding
         --         to the real space resolution <R3d>.
    ---C++: inline
    ;   
        
    GetType(myclass; C: HCurve2d from Adaptor2d) returns CurveType from GeomAbs
	---Purpose: Returns  the  type of the   curve  in the  current
	--          interval :   Line,   Circle,   Ellipse, Hyperbola,
	--          Parabola, BezierCurve, BSplineCurve, OtherCurve.
    ---C++: inline
    ;

    --
    --     The following methods must  be called when GetType returned
    --     the corresponding type.
    --     

     Line(myclass; C: HCurve2d from Adaptor2d) returns Lin2d from gp
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;
     
     Circle(myclass; C: HCurve2d from Adaptor2d) returns Circ2d from gp
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;
     
     Ellipse(myclass; C: HCurve2d from Adaptor2d) returns Elips2d from gp
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;
     
     Hyperbola(myclass; C: HCurve2d from Adaptor2d) returns  Hypr2d from gp
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;
     
     Parabola(myclass; C: HCurve2d from Adaptor2d) returns Parab2d from gp
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;
     
     Bezier(myclass; C: HCurve2d from Adaptor2d) returns BezierCurve from Geom2d
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;
    
     BSpline(myclass; C: HCurve2d from Adaptor2d) returns BSplineCurve from Geom2d
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;

    



    NbSamples(myclass; C: HCurve2d from Adaptor2d; U0,U1: Real from Standard) 
    returns Integer from Standard;

end HCurve2dTool;
