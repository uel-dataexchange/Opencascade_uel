-- File:        SeamCurve.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSeamCurve from RWStepGeom

	---Purpose : Read & Write Module for SeamCurve

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SeamCurve from StepGeom,
     EntityIterator from Interface

is

	Create returns RWSeamCurve;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable SeamCurve from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : SeamCurve from StepGeom);

	Share(me; ent : SeamCurve from StepGeom; iter : in out EntityIterator);

end RWSeamCurve;
