-- File:	StepToGeom_MakeDirection.cdl
-- Created:	Mon Jun 14 14:53:21 1993
-- Author:	Martine LANGLOIS
---Copyright:	 Matra Datavision 1993

class MakeDirection from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          Direction from StepGeom which describes a direction
    --          from Prostep and Direction from Geom.

uses 
     Direction from Geom,
     Direction from StepGeom

is 

    Convert ( myclass; SD : Direction from StepGeom;
                       CD : out Direction from Geom )
    returns Boolean from Standard;

end MakeDirection;
