-- File:	RWStepBasic_RWConversionBasedUnitAndVolumeUnit.cdl
-- Created:	Tue Oct 12 14:28:52 1999
-- Author:	data exchange team
--		<det@friendox>
---Copyright:	 Matra Datavision 1999


class RWConversionBasedUnitAndVolumeUnit from RWStepBasic 

	---Purpose: Read & Write Module for ConversionBasedUnitAndVolumeUnit

uses

    Check from Interface,
    StepReaderData from StepData,
    StepWriter from StepData,
    ConversionBasedUnitAndVolumeUnit from StepBasic,
    EntityIterator from Interface

is

    Create returns RWConversionBasedUnitAndVolumeUnit from RWStepBasic;
    
    ReadStep (me; data: StepReaderData; num : Integer;
	          ach : in out Check; ent : mutable ConversionBasedUnitAndVolumeUnit from StepBasic);

    WriteStep (me; SW : in out StepWriter; ent : ConversionBasedUnitAndVolumeUnit from StepBasic);

    Share(me; ent : ConversionBasedUnitAndVolumeUnit from StepBasic; iter : in out EntityIterator);


end RWConversionBasedUnitAndVolumeUnit;
