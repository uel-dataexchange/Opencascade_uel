-- File:        PresentationSet.cdl
-- Created:     Fri Dec  1 11:11:25 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class PresentationSet from StepVisual 

inherits TShared from MMgt

is

	Create returns mutable PresentationSet;
	---Purpose: Returns a PresentationSet


end PresentationSet;
