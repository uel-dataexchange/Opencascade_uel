-- File:	RWStepAP214_RWAppliedApprovalAssignment.cdl
-- Created:	Fri Mar 12 11:44:44 1999
-- Author:	data exchange team
--		<det@androx.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class RWAppliedApprovalAssignment from RWStepAP214 

	---Purpose: Read & Write Module for AppliedApprovalAssignment

uses
     Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     AppliedApprovalAssignment from StepAP214,
     EntityIterator from Interface


is
    	Create returns RWAppliedApprovalAssignment;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable AppliedApprovalAssignment from StepAP214);

	WriteStep (me; SW : in out StepWriter; ent : AppliedApprovalAssignment from StepAP214);

	Share(me; ent : AppliedApprovalAssignment from StepAP214; iter : in out EntityIterator);


end RWAppliedApprovalAssignment;
