-- File:	FairCurve_EnergyOfMVC.cdl
-- Created:	Mon Apr  1 09:10:45 1996
-- Author:	Philippe MANGIN
--		<pmn@sgi29>
---Copyright:	 Matra Datavision 1996


private class EnergyOfMVC from FairCurve  inherits Energy from FairCurve

	---Purpose: Energy Criterium to minimize in MinimalVariationCurve.
	---Category: Private use

uses BattenLaw from FairCurve,  
     DistributionOfTension from FairCurve, 
     DistributionOfSagging from FairCurve,
     DistributionOfJerk    from FairCurve,
     AnalysisCode from FairCurve,
     Vector  from  math,
     Matrix  from math,
     HArray1OfPnt2d from TColgp,
     Array1OfXY  from TColgp,
     Pnt2d from gp,
     HArray1OfReal from TColStd
     
raises DomainError


is
    Create( BSplOrder     : Integer;
            FlatKnots     : HArray1OfReal;
	    Poles         : HArray1OfPnt2d;
    	    ContrOrder1   : Integer;
	    ContrOrder2   : Integer;
	    Law           : BattenLaw;
	    PhysicalRatio : Real;
	    LengthSliding : Real;
	    FreeSliding   : Boolean = Standard_True;
            Angle1        : Real = 0;
            Angle2        : Real = 0;
    	    Curvature1    : Real = 0;
    	    Curvature2    : Real = 0 )
     ---Purpose: Angles corresspond to the Ox axis
     returns  EnergyOfMVC
     raises  DomainError; -- if  PhysicalRatio < 0 or  PhysicalRatio > 1
    
    LengthSliding(me)
    ---Purpose: return  the  lengthSliding = P1P2 + Sliding
    ---C++: inline
    returns  Real;
    
         
    Status(me) 
    ---Purpose: return  the status 
    ---C++: inline
    returns  AnalysisCode;
    
    ComputePoles(me: in out; X: Vector)
    ---Purpose: compute  the  poles wich correspond with the variable X
    is redefined protected; 
    
    Variable(me; X: out Vector)
    ---Purpose: compute the variables <X> wich correspond with the field <MyPoles>
    returns Boolean
    is redefined;  
	
    Compute(me:in out; DerivativeOrder : Integer; Result : out Vector)
        ---Purpose: compute the energy in intermediat format
    returns Boolean 
    is redefined protected;
    
fields
    MyLengthSliding : Real;
    OriginalSliding : Real;
    MyFreeSliding   : Boolean;
    MyBattenLaw     : BattenLaw;
    MyPhysicalRatio : Real;
    MyTension       : DistributionOfTension;
    MySagging       : DistributionOfSagging;
    MyJerk          : DistributionOfJerk;
    MyStatus        : AnalysisCode;

end EnergyOfMVC;
