-- File:	RWStepShape_RWDimensionalLocationWithPath.cdl
-- Created:	Tue Apr 18 16:42:58 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWDimensionalLocationWithPath from RWStepShape

    ---Purpose: Read & Write tool for DimensionalLocationWithPath

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    DimensionalLocationWithPath from StepShape

is
    Create returns RWDimensionalLocationWithPath from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : DimensionalLocationWithPath from StepShape);
	---Purpose: Reads DimensionalLocationWithPath

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: DimensionalLocationWithPath from StepShape);
	---Purpose: Writes DimensionalLocationWithPath

    Share (me; ent : DimensionalLocationWithPath from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWDimensionalLocationWithPath;
