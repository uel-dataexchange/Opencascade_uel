-- File:      XmlMFunction_ScopeDriver.cdl
-- Created:   04.03.08 15:37:51
-- Author:    Vlad ROMASHKO
-- Copyright: Open Cascade 2008

class ScopeDriver from XmlMFunction  inherits ADriver from XmlMDF

        ---Purpose: XML persistence driver for a scope of functions.

uses

    SRelocationTable from XmlObjMgt,
    RRelocationTable from XmlObjMgt,
    Persistent       from XmlObjMgt,
    MessageDriver    from CDM,
    Attribute        from TDF

is

    Create (theMessageDriver : MessageDriver from CDM)
    returns mutable ScopeDriver from XmlMFunction;

    NewEmpty (me)  
    returns mutable Attribute from TDF;

    Paste(me; Source     : Persistent from XmlObjMgt;
              Target     : mutable Attribute from TDF;
              RelocTable : out RRelocationTable from XmlObjMgt)
    returns Boolean from Standard;

    Paste(me; Source     : Attribute from TDF;
              Target     : in out Persistent from XmlObjMgt;
              RelocTable : out SRelocationTable from XmlObjMgt);

end ScopeDriver;
