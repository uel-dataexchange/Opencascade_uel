-- File:	STEPCAFControl_Writer.cdl
-- Created:	Tue Aug 15 17:23:00 2000
-- Author:	Andrey BETENEV
--		<abv@doomox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2000


class Writer from STEPCAFControl 
-- inherits Writer from STEPControl

    ---Purpose: Provides a tool to write DECAF document to the
    --          STEP file. Besides transfer of shapes (including 
    --          assemblies) provided by STEPControl, supports also 
    --          colors and part names
    --
    --          Also supports multifile writing

uses
    AsciiString from TCollection,
    ReturnStatus from IFSelect,
    WorkSession from XSControl,
    Shape from TopoDS,
    Writer from STEPControl,
    StepModelType from STEPControl,
    DictionaryOfExternFile from STEPCAFControl,
    ExternFile from STEPCAFControl,
    Label from TDF,
    LabelSequence from TDF,
    DataMapOfLabelShape from STEPCAFControl,
    DataMapOfLabelExternFile from STEPCAFControl,
    Document from TDocStd,
    DataMapOfShapeTransient from MoniTool

is

    Create returns Writer;
    	---Purpose: Creates a writer with an empty
-- STEP model and sets ColorMode, LayerMode, NameMode and
-- PropsMode to Standard_True.
        
    Create (WS : mutable WorkSession from XSControl;
    	    	 scratch : Boolean = Standard_True) returns Writer;
    	---Purpose: Creates a reader tool and attaches it to an already existing Session
    	--          Clears the session if it was not yet set for STEP
	--          Clears the internal data structures

    Init (me: in out; WS : mutable WorkSession from XSControl;
    	              scratch : Boolean = Standard_True);
    	---Purpose: Clears the internal data structures and attaches to a new session
    	--          Clears the session if it was not yet set for STEP

    Write (me : in out; filename : CString) 
    returns ReturnStatus from IFSelect;
        ---Purpose: Writes all the produced models into file
	--          In case of multimodel with extern references,
	--          filename will be a name of root file, all other files
	--          have names of corresponding parts
	--          Provided for use like single-file writer

    Transfer (me : in out; doc : Document from TDocStd;
    	    	    	   mode: StepModelType from STEPControl = STEPControl_AsIs;
			   multi: CString = 0)
    returns Boolean;
    Transfer (me : in out; L: Label from TDF;
    	    	    	   mode: StepModelType from STEPControl = STEPControl_AsIs;
			   multi: CString = 0)
    returns Boolean;
    	---Purpose: Transfers a document (or single label) to a STEP model
    	--          The mode of translation of shape is AsIs
	--          If multi is not null pointer, it switches to multifile
	--          mode (with external refs), and string pointed by <multi>
	--          gives prefix for names of extern files (can be empty string)
    	--          Returns True if translation is OK

    Perform (me : in out; doc : Document from TDocStd;
    	    	    	  filename: AsciiString from TCollection)
    returns Boolean;

    Perform (me : in out; doc : Document from TDocStd; filename: CString)
    returns Boolean;
    ---Purpose : Transfers a document and writes it to a STEP file
    --           Returns True if translation is OK

    ---Scope: Access to fields
    
    ExternFiles (me) returns DictionaryOfExternFile from STEPCAFControl;
    	---Purpose: Returns data on external files
	--          Returns Null handle if no external files are read
	---C++: return const &
	
    ExternFile (me; L: Label from TDF; ef: out ExternFile from STEPCAFControl)
    returns Boolean;
    	---Purpose: Returns data on external file by its original label
	--          Returns False if no external file with given name is read
	
    ExternFile (me; name: CString; ef: out ExternFile from STEPCAFControl)
    returns Boolean;
    	---Purpose: Returns data on external file by its name
	--          Returns False if no external file with given name is read
	
    ChangeWriter (me: in out) returns Writer from STEPControl;
    	---Purpose: Returns basic reader for root file
	---C++: return &

    Writer (me) returns Writer from STEPControl;
    	---Purpose: Returns basic reader as const
	---C++: return const &

    ---Scope: Internal methods

    Transfer (me : in out; wr: in out Writer from STEPControl;
    	    	    	   labels: LabelSequence from TDF;
    	    	    	   mode: StepModelType from STEPControl = STEPControl_AsIs;
			   multi: CString = 0;
    	    	    	   isExternFile: Boolean = Standard_False)
    returns Boolean is protected;
    	---Purpose: Transfers labels to a STEP model
    	--          Returns True if translation is OK
	--          isExternFile setting from TransferExternFiles method

    TransferExternFiles (me : in out; L: Label from TDF;
    	    	    	              mode: StepModelType from STEPControl;
			              Lseq: out LabelSequence from TDF;
    	    	    	    	      prefix: CString = "")
    returns Shape from TopoDS is protected;
    	---Purpose: Parses assembly structure of label L, writes all the simple
        --          shapes each to its own file named by name of its label plus
        --          prefix
        --          Returns shape representing that assembly structure
        --          in the form of nested empty compounds (and a sequence of 
	--          labels which are newly written nodes of this assembly)

    WriteExternRefs (me; WS: WorkSession from XSControl; labels: LabelSequence from TDF) 
    returns Boolean is protected;
    	---Purpose: Write external references to STEP

    WriteColors (me: in out; WS: WorkSession from XSControl; labels: LabelSequence from TDF) 
    returns Boolean is protected;
    	---Purpose: Write colors assigned to specified labels, to STEP model

    WriteNames (me; WS: WorkSession from XSControl; labels: LabelSequence from TDF) 
    returns Boolean is protected;
    	---Purpose: Write names assigned to specified labels, to STEP model

    WriteDGTs (me; WS: WorkSession from XSControl; labels: LabelSequence from TDF) 
    returns Boolean is protected;
    	---Purpose: Write D&GTs assigned to specified labels, to STEP model

    WriteMaterials (me; WS: WorkSession from XSControl; labels: LabelSequence from TDF) 
    returns Boolean is protected;
    	---Purpose: Write materials assigned to specified labels, to STEP model

    WriteValProps (me; WS: WorkSession from XSControl; 
                       labels: LabelSequence from TDF; multi: CString)
    returns Boolean is protected;
    	---Purpose: Write validation properties assigned to specified labels, 
        --          to STEP model

    WriteLayers (me; WS: WorkSession from XSControl; labels: LabelSequence from TDF) 
    returns Boolean is protected;
    	---Purpose: Write layers assigned to specified labels, to STEP model

    WriteSHUOs (me: in out; WS: WorkSession from XSControl; labels: LabelSequence from TDF)
    returns Boolean is protected;
    	---Purpose: Write SHUO assigned to specified component, to STEP model

    --- Work with fileds for different mode of writing STEP file.

    SetColorMode(me: in out; colormode: Boolean from Standard);
    	---Purpose: Set ColorMode for indicate write Colors or not.

    GetColorMode(me) returns Boolean;

    SetNameMode(me: in out; namemode: Boolean from Standard);
    	---Purpose: Set NameMode for indicate write Name or not.
    
    GetNameMode(me) returns Boolean;

    SetLayerMode(me: in out; layermode: Boolean from Standard);
    	---Purpose: Set LayerMode for indicate write Layers or not.

    GetLayerMode(me) returns Boolean; 
    
    SetPropsMode(me: in out; propsmode: Boolean from Standard);
    	---Purpose: PropsMode for indicate write Validation properties or not.

    GetPropsMode(me) returns Boolean;
	
    SetSHUOMode(me: in out; shuomode: Boolean from Standard);
    	---Purpose: Set SHUO mode for indicate write SHUO or not.

    GetSHUOMode(me) returns Boolean;
	
    SetDimTolMode(me: in out; dimtolmode: Boolean from Standard);
    	---Purpose: Set dimtolmode for indicate write D&GTs or not.

    GetDimTolMode(me) returns Boolean;
	
    SetMaterialMode(me: in out; matmode: Boolean from Standard);
    	---Purpose: Set dimtolmode for indicate write D&GTs or not.

    GetMaterialMode(me) returns Boolean;
	
fields

    myWriter : Writer from STEPControl;
    myFiles  : DictionaryOfExternFile from STEPCAFControl;
    myLabels : DataMapOfLabelShape from STEPCAFControl;
    myLabEF  : DataMapOfLabelExternFile from STEPCAFControl;
    myColorMode: Boolean;
    myNameMode : Boolean;
    myLayerMode: Boolean;
    myPropsMode: Boolean;
    mySHUOMode : Boolean;
    myMapCompMDGPR : DataMapOfShapeTransient from MoniTool;
    myDGTMode  : Boolean;
    myMatMode  : Boolean;

end Writer;
