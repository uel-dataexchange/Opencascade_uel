--
-- File:	AlienImage_EuclidAlienImage.cdl
-- Created:	23/03/93
-- Author:	BBL
-- Modified:	02-06-98 : FMN ; Suppression appel Clear (deja fait dans ALienData)
--
---Copyright:	Matravision 1993
--

class EuclidAlienImage from AlienImage inherits AlienUserImage from AlienImage

	---Version: 0.0

	---Purpose: This class defines an Euclid Alien image.
	---Keywords:
	---Warning:
	---References:

uses
	File 			from OSD,
	AsciiString 		from TCollection,
	ColorImage 		from Image,
	PseudoColorImage 	from Image,
	Image			from Image,
	EuclidAlienData 	from AlienImage

is
	Create returns mutable EuclidAlienImage from AlienImage;

	Clear( me : in out mutable) ;
	---Level: Public
	---Purpose: Frees memory allocated by EuclidAlienImage

	ToImage( me : in immutable ) 
	  returns mutable Image from Image ;
	---Level: Public
	---Purpose : Converts a EuclidAlienImage object to a Image object.

	FromImage( me : in out mutable ; anImage : in Image from Image ) ;
	---Level: Public
	---Purpose : converts a Image object to a EuclidAlienImage object.

	Read ( me : in out mutable; afile : in out File from OSD )
	  returns Boolean from Standard ;
	---Purpose: Reads content of a EuclidAlienImage object
	--          from a file .
	--          Returns True if file is a Euclid file .

	Write( me : in immutable; afile : in out File from OSD )
	  returns Boolean from Standard ;
	---Purpose: Writes content of a EuclidAlienImage object
	--          to a file .

fields
	myData : EuclidAlienData from AlienImage ;

end ;
 
