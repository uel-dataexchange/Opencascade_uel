-- File:	BOP_LoopClassifier.cdl
-- Created:	Wed Mar  3 17:29:13 1993
-- Author:	Jean Yves LEBEY
--		<jyl@sdsun2>
---Copyright:	 Matra Datavision 1993

deferred class LoopClassifier from BOP 

    ---Purpose:  
    --  Root class to classify Loops in order to build Areas

uses

    ShapeEnum from TopAbs,
    State from TopAbs,
    Loop from BOP
    
is

    Delete(me:out) is virtual;
    	---C++: alias "Standard_EXPORT virtual ~BOP_LoopClassifier(){Delete() ; }"
    	---Purpose:  
    	--- Destructor;  
    	---
    Compare(me : in out; L1,L2 : Loop from BOP) 
    	returns State from TopAbs  
    	is deferred;
    	---Purpose:  
    	--- Returns the state of loop <L1> compared with loop <L2>.
    	---
    
end LoopClassifier;
