-- File:        PresentationView.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPresentationView from RWStepVisual

	---Purpose : Read & Write Module for PresentationView

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PresentationView from StepVisual,
     EntityIterator from Interface

is

	Create returns RWPresentationView;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PresentationView from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : PresentationView from StepVisual);

	Share(me; ent : PresentationView from StepVisual; iter : in out EntityIterator);

end RWPresentationView;
