-- File:        FaceBound.cdl
-- Created:     Mon Dec  4 12:02:26 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWFaceBound from RWStepShape

	---Purpose : Read & Write Module for FaceBound
	--           Check added by CKY , 7-OCT-1996

uses Check from Interface, ShareTool from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     FaceBound from StepShape,
     EntityIterator from Interface

is

	Create returns RWFaceBound;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable FaceBound from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : FaceBound from StepShape);

	Share(me; ent : FaceBound from StepShape; iter : in out EntityIterator);

	Check(me; ent : FaceBound from StepShape; shares : ShareTool; ach : in out Check);

end RWFaceBound;
