-- File:	Dynamic_BooleanParameter.cdl
-- Created:	Mon Jan 24 13:33:06 1994
-- Author:	Gilles DEBARBOUILLE
--		<gde@meteox>
---Copyright:	 Matra Datavision 1994


class BooleanParameter from Dynamic

inherits
    Parameter from Dynamic     
    
	---Purpose: This class describes a parameter with a boolean 
	--          as value.

uses

   CString from Standard,
   OStream from Standard

is

    Create(aparameter : CString from Standard)
    
    ---Level: Advanced 
    
    ---Purpose: Creates a boolean parameter with <aparameter> as name.

    returns mutable BooleanParameter from Dynamic;
    
    Create(aparameter : CString from Standard; 
           avalue : Boolean from Standard) 

    ---Level: Advanced 
    
    ---Purpose: Creates a boolean parameter with <aparameter> and <avalue>
    --          respectively as name and value.

    returns mutable BooleanParameter from Dynamic;
    
    Create(aparameter , avalue : CString from Standard)
    
    ---Level: Advanced 
    
    ---Purpose: Creates a boolean parameter with <aparameter> as name 
    --          and <avalue> as value. <avalue> is a CString with two possible
    --          values which are : "Standard_True" and "Standard_False".

    returns mutable BooleanParameter from Dynamic;
    
    Value(me) returns Boolean from Standard
    
    ---Level: Public 
    
    ---Purpose: Returns the boolean value <thevalue>.
    
    is static;
    
    Value (me : mutable ; avalue : Boolean from Standard)
    
    ---Level: Advanced 
    
    --- Purpose: Sets the field <thevalue> with the boolean value <avalue>

    is static;
    
    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Internal 
    
    ---Purpose: Useful for debugging.
    
    is redefined;
    
fields

    thevalue : Boolean from Standard;

end BooleanParameter;
