-- File:	StepRepr_DataEnvironment.cdl
-- Created:	Thu Dec 12 15:38:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class DataEnvironment from StepRepr
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity DataEnvironment

uses
    HAsciiString from TCollection,
    HArray1OfPropertyDefinitionRepresentation from StepRepr

is
    Create returns DataEnvironment from StepRepr;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       aDescription: HAsciiString from TCollection;
                       aElements: HArray1OfPropertyDefinitionRepresentation from StepRepr);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

    Elements (me) returns HArray1OfPropertyDefinitionRepresentation from StepRepr;
	---Purpose: Returns field Elements
    SetElements (me: mutable; Elements: HArray1OfPropertyDefinitionRepresentation from StepRepr);
	---Purpose: Set field Elements

fields
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection;
    theElements: HArray1OfPropertyDefinitionRepresentation from StepRepr;

end DataEnvironment;
