-- File:        CoordinatedUniversalTimeOffset.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWCoordinatedUniversalTimeOffset from RWStepBasic

	---Purpose : Read & Write Module for CoordinatedUniversalTimeOffset

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     CoordinatedUniversalTimeOffset from StepBasic

is

	Create returns RWCoordinatedUniversalTimeOffset;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable CoordinatedUniversalTimeOffset from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : CoordinatedUniversalTimeOffset from StepBasic);

end RWCoordinatedUniversalTimeOffset;
