-- File:        PointReplica.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPointReplica from RWStepGeom

	---Purpose : Read & Write Module for PointReplica

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PointReplica from StepGeom,
     EntityIterator from Interface

is

	Create returns RWPointReplica;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PointReplica from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : PointReplica from StepGeom);

	Share(me; ent : PointReplica from StepGeom; iter : in out EntityIterator);

end RWPointReplica;
