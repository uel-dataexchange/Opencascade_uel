-- File:	RWStepBasic_RWExternallyDefinedItem.cdl
-- Created:	Wed May 10 15:09:07 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWExternallyDefinedItem from RWStepBasic

    ---Purpose: Read & Write tool for ExternallyDefinedItem

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ExternallyDefinedItem from StepBasic

is
    Create returns RWExternallyDefinedItem from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ExternallyDefinedItem from StepBasic);
	---Purpose: Reads ExternallyDefinedItem

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ExternallyDefinedItem from StepBasic);
	---Purpose: Writes ExternallyDefinedItem

    Share (me; ent : ExternallyDefinedItem from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWExternallyDefinedItem;
