-- File:	MXCAFDoc_DimTolStorageDriver.cdl
-- Created:	Wed Dec 10 09:05:14 2008
-- Author:	Pavel TELKOV
--		<ptv@valenox>
---Copyright:	 Open CASCADE 2008

class DimTolStorageDriver from MXCAFDoc inherits ASDriver from MDF

	---Purpose: 
uses
    SRelocationTable from MDF,
    Attribute        from TDF,
    Attribute        from PDF,
    MessageDriver    from CDM

is

    Create (theMsgDriver : MessageDriver from CDM)
    returns mutable DimTolStorageDriver from MXCAFDoc;
	---Purpose: Returns mutable DimTolStorageDriver from MXCAFDoc;

    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type: XCAFDoc_DimTol.

    NewEmpty (me) returns mutable Attribute from PDF;

    Paste(me;
    	  Source     :         Attribute from TDF;
    	  Target     : mutable Attribute from PDF;
    	  RelocTable : SRelocationTable from MDF);

end DimTolStorageDriver;
