-- File:	RWStepFEA_RWElementGroup.cdl
-- Created:	Thu Dec 12 17:51:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWElementGroup from RWStepFEA

    ---Purpose: Read & Write tool for ElementGroup

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ElementGroup from StepFEA

is
    Create returns RWElementGroup from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ElementGroup from StepFEA);
	---Purpose: Reads ElementGroup

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ElementGroup from StepFEA);
	---Purpose: Writes ElementGroup

    Share (me; ent : ElementGroup from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWElementGroup;
