-- File:        LimitsAndFits.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWLimitsAndFits from RWStepShape

	---Purpose : Read & Write Module for LimitsAndFits

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     LimitsAndFits from StepShape

is

	Create returns RWLimitsAndFits;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable LimitsAndFits from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : LimitsAndFits from StepShape);

end RWLimitsAndFits;
