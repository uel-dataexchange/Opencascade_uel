-- File:	RWStepBasic_RWExternalIdentificationAssignment.cdl
-- Created:	Wed May 10 15:09:06 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWExternalIdentificationAssignment from RWStepBasic

    ---Purpose: Read & Write tool for ExternalIdentificationAssignment

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ExternalIdentificationAssignment from StepBasic

is
    Create returns RWExternalIdentificationAssignment from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ExternalIdentificationAssignment from StepBasic);
	---Purpose: Reads ExternalIdentificationAssignment

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ExternalIdentificationAssignment from StepBasic);
	---Purpose: Writes ExternalIdentificationAssignment

    Share (me; ent : ExternalIdentificationAssignment from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWExternalIdentificationAssignment;
