-- File:        SurfaceStyleBoundary.cdl
-- Created:     Fri Dec  1 11:11:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class SurfaceStyleBoundary from StepVisual 

inherits TShared from MMgt

uses

	CurveStyle from StepVisual
is

	Create returns mutable SurfaceStyleBoundary;
	---Purpose: Returns a SurfaceStyleBoundary

	Init (me : mutable;
	      aStyleOfBoundary : mutable CurveStyle from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetStyleOfBoundary(me : mutable; aStyleOfBoundary : mutable CurveStyle);
	StyleOfBoundary (me) returns mutable CurveStyle;

fields

	styleOfBoundary : CurveStyle from StepVisual;

end SurfaceStyleBoundary;
