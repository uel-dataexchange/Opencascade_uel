-- File:        DraughtingPreDefinedColour.cdl
-- Created:     Fri Dec  1 11:11:19 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class DraughtingPreDefinedColour from StepVisual 

inherits PreDefinedColour from StepVisual 

uses

	HAsciiString from TCollection
is

	Create returns mutable DraughtingPreDefinedColour;
	---Purpose: Returns a DraughtingPreDefinedColour


end DraughtingPreDefinedColour;
