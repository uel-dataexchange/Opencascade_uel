-- File:	NLPlate_HPG0G3Constraint.cdl
-- Created:	Fri Apr 17 15:11:16 1998
-- Author:	Andre LIEUTIER
--		<alr@sgi63>
---Copyright:	 Matra Datavision 1998



class  HPG0G3Constraint  from  NLPlate  inherits  HPG0G2Constraint from  NLPlate 
---Purpose: define a PinPoint G0+G3  Constraint  used to load a Non Linear
--          Plate
uses
     XY from gp,
     XYZ from gp, 
     D1  from  Plate,
     D2  from  Plate,
     D3  from  Plate
     
is
    Create(UV : XY; Value : XYZ; D1T : D1 from Plate; 
     D2T : D2 from Plate;  D3T : D3 from Plate) returns mutable HPG0G3Constraint;
    -- create a G0+G3 Constraint
    -- 

    ActiveOrder(me)  returns  Integer 
    is   redefined; 
    --  returns the constraint active  order, i.e. the maximum between
    --  -- the initial constraint i.e 3 (for G3 Constraints)

 
    G3Target(me) returns D3 from Plate
    ---C++: return const &
    is  redefined; 
        

fields
     myG3Target : D3 from Plate; 
end;
