-- File:	GProp_FaceTool.cdl
-- Created:	Fri Nov 27 16:29:37 1992
-- Author:	Isabelle GRIGNON
--		<isg@sdsun2>
---Copyright:	 Matra Datavision 1992

deferred generic class FaceTool  from GProp( Arc as any )

        ---Purpose: This template class defines the minimum of methods required 
        --          to compute the global properties of Faces with the 
        --          algorithms of the package GProp. 
        --          To compute the global properties of a Face, in is necessary
        --          to define own "FaceTool" and to implement all the methods 
        --          defined in this template. Note that it is not necessary to 
        --          inherit this template class.
	
uses Pnt           from gp,
     Pnt2d         from gp,
     Vec           from gp,
     Vec2d         from gp, 
     IsoType       from GeomAbs, 
     HArray1OfReal from TColStd

is 

  UIntegrationOrder (me) returns Integer;
        ---Purpose: Returns the number of points required to do the 
        --          integration in the U parametric direction.

  Bounds (me; U1, U2, V1, V2 : out Real);
	---Purpose: Returns the parametric bounds of the Face <S>.

  Normal (me;  U, V : Real; P : out Pnt; VNor: out Vec);
	---Purpose: Computes the point of parameter U, V on the Face <S> and 
	--          the normal to the face at this point.

  Load(me:in out; A : Arc); 
        ---Purpose: Loading the boundary arc.
  
  Load(me : in out; IsFirstParam: Boolean from Standard; 
                    theIsoType  : IsoType from GeomAbs);
        ---Purpose: Loading the boundary arc. This arc is either a top, bottom, 
        --          left or right bound of a UV rectangle in which the 
        --          parameters of surface are defined. 
	--          If IsFirstParam is equal to Standard_True, the face is 
        --          initialized by either left of bottom bound. Otherwise it is 
        --          initialized by the top or right one. 
	--          If theIsoType is equal to GeomAbs_IsoU, the face is 
        --          initialized with either left or right bound. Otherwise - 
        --          with either top or bottom one.
  
  FirstParameter (me) returns Real ;
        ---Purpose: Returns the parametric value of the start point of
        --          the current arc of curve. 

  LastParameter (me) returns Real ;
        ---Purpose: Returns the parametric value of the end point of
        --          the current arc of curve. 

  IntegrationOrder (me) returns Integer;
        ---Purpose: Returns the number of points required to do the 
        --          integration along the parameter of curve.

  D12d (me; U: Real; P: out Pnt2d; V1: out Vec2d);
    	---Purpose: Returns the point of parameter U and the first derivative 
    	--          at this point of a boundary curve.

  GetUKnots(me; theUMin  :        Real          from Standard; 
                theUMax  :        Real          from Standard; 
		theUKnots: in out HArray1OfReal from TColStd); 
	---Purpose: Returns an array of U knots of the face. The first and last 
        --          elements of the array will be theUMin and theUMax. The 
        --          middle elements will be the U Knots of the face greater 
        --          then theUMin and lower then theUMax in increasing order. 

  GetTKnots(me; theTMin  :        Real          from Standard; 
                theTMax  :        Real          from Standard; 
		theTKnots: in out HArray1OfReal from TColStd);
	---Purpose: Returns an array of combination of T knots of the arc and 
        --          V knots of the face. The first and last elements of the 
        --          array will be theTMin and theTMax. The middle elements will 
        --          be the Knots of the arc and the values of parameters of 
        --          arc on which the value points have V coordinates close to V 
        --          knots of face. All the parameter will be greater then 
        --          theTMin and lower then theTMax in increasing order.

end FaceTool;









