-- File:	StepElement_Surface3dElementDescriptor.cdl
-- Created:	Thu Dec 12 17:29:04 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class Surface3dElementDescriptor from StepElement
inherits ElementDescriptor from StepElement

    ---Purpose: Representation of STEP entity Surface3dElementDescriptor

uses
    ElementOrder from StepElement,
    HAsciiString from TCollection,
    HArray1OfHSequenceOfSurfaceElementPurposeMember from StepElement,
    Element2dShape from StepElement

is
    Create returns Surface3dElementDescriptor from StepElement;
	---Purpose: Empty constructor

    Init (me: mutable; aElementDescriptor_TopologyOrder: ElementOrder from StepElement;
                       aElementDescriptor_Description: HAsciiString from TCollection;
                       aPurpose: HArray1OfHSequenceOfSurfaceElementPurposeMember from StepElement;
                       aShape: Element2dShape from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    Purpose (me) returns HArray1OfHSequenceOfSurfaceElementPurposeMember from StepElement;
	---Purpose: Returns field Purpose
    SetPurpose (me: mutable; Purpose: HArray1OfHSequenceOfSurfaceElementPurposeMember from StepElement);
	---Purpose: Set field Purpose

    Shape (me) returns Element2dShape from StepElement;
	---Purpose: Returns field Shape
    SetShape (me: mutable; Shape: Element2dShape from StepElement);
	---Purpose: Set field Shape

fields
    thePurpose: HArray1OfHSequenceOfSurfaceElementPurposeMember from StepElement;
    theShape: Element2dShape from StepElement;

end Surface3dElementDescriptor;
