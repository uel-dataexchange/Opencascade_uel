-- File:	Dynamic_CompiledMethod.cdl
-- Created:	Thu Jan 28 14:59:01 1993
-- Author:	Gilles DEBARBOUILLE
--		<gde@bravox>
---Copyright:	 Matra Datavision 1993


class CompiledMethod from Dynamic

inherits

    MethodDefinition from Dynamic
    ---Purpose: A Dynamic_CompiledMethod adds to the definition of the
    --          Dynamic_Method the C++ mangled name of the function to
    --          be  run. An application using  instances of this class
    --          must bind the C++  name of  the  method with the  true
    --          address in the executable.

uses

    CString from Standard,
    HAsciiString from TCollection,
    AsciiString  from TCollection


is

    Create(aname : CString from Standard;
           afunction : CString from Standard) returns mutable CompiledMethod from Dynamic;
    
    ---Level: Advanced 
    
    ---Purpose: Creates  a compiled method   with <aname> as user name
    --          and <afunction> as C++ mangled name.
    
    Function(me : mutable ; afunction : CString from Standard)
    
    ---Level: Advanced 
    
    ---Purpose: Sets the  C++ mangled name  of the method to the field
    --          <thefunction>.
    
    is static;
    
    Function(me) returns AsciiString from TCollection
    
    ---Level: Advanced 
    
    ---Purpose: Returns the C++ mangled name of the function.
    
    is static;
    
fields

    thefunction : HAsciiString from TCollection;

end CompiledMethod;
