-- File:	IGESSelect_SelectFromSingleView.cdl
-- Created:	Tue May 31 18:36:13 1994
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1994


class SelectFromSingleView  from IGESSelect  inherits SelectDeduct

    ---Purpose : This selection gets in all the model, the entities which are
    --           attached to the views given as input. Only Single Views are
    --           considered. This information is kept from Directory Part
    --           (View Item).

uses AsciiString from TCollection, EntityIterator, Graph

raises InterfaceError

is

    Create returns mutable SelectFromSingleView;
    ---Purpose : Creates a SelectFromSingleView

    RootResult (me; G : Graph) returns EntityIterator  raises InterfaceError;
    ---Purpose : Selects the Entities which are attached to the Single View(s)
    --           present in the Input

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns the label, with is "Entities attached to single View"

end SelectFromSingleView;
