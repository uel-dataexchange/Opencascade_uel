-- File:      BRepExtrema.cdl
-- Created:   Fri Dec  3 15:48:19 1993
-- Author:    Christophe MARION
---Copyright: Matra Datavision 1993

package BRepExtrema

    ---Purpose: This package gives   tools to compute  extrema between
    --          Shapes from BRep.

uses 
    Standard,
    StdFail,
    TopoDS,
    GeomAdaptor,
    BRepAdaptor,
    gp,
    Extrema,
    TColStd,
    TopTools,
    TCollection,
    Bnd
    
is

    ----------------------------------------------------------
    --  Extrema between two Shapes with triangulation.
    ----------------------------------------------------------
    imported Poly;


    ----------------------------------------------------------
    --  Extrema between a Point and an Edge.
    ----------------------------------------------------------
    imported ExtPC;


    ----------------------------------------------------------
    --  Extrema between two Edges.
    ----------------------------------------------------------
    imported ExtCC;


    ----------------------------------------------------------
    --  Extrema between a Point and a Face.
    ----------------------------------------------------------
    imported ExtPF;


    ----------------------------------------------------------
    --  Extrema between an Edge  and a Face.
    ----------------------------------------------------------
    imported ExtCF;


    ----------------------------------------------------------
    --  Extrema between two Faces.
    ----------------------------------------------------------
    imported ExtFF;


    ----------------------------------------------------------
    --  
    ----------------------------------------------------------
    exception UnCompatibleShape inherits DomainError;


    ----------------------------------------------------------
    --  enumeration used to describe the type of the support solution:                                         
    -- 	    IsVertex => The solution is a vertex.
    -- 	    IsOnEdge => The solution belongs to an Edge.
    -- 	    IsInFace => The solution is inside a Face.    
     
    ----------------------------------------------------------
    imported SupportType;


    ----------------------------------------------------------
    -- This  class gives tools  to  compute the minimum distance value
    -- between two shapes and  the corresponding couples of solution points.  
    
    ----------------------------------------------------------
    imported DistShapeShape;


    ----------------------------------------------------------
    --  This class is used to store a solution on a Shape. 
    --  (used only by class DistShapeShape)
    ----------------------------------------------------------
    imported SolutionElem;


    ----------------------------------------------------------
    -- This sequence is used to store all the solution on each Shape.
    ----------------------------------------------------------
    imported SeqOfSolution;

    imported DistanceSS;

end BRepExtrema;
