-- File:	MDataStd_AsciiStringRetrievalDriver.cdl
-- Created:	Thu Aug 23 09:55:00 2007
-- Author:	Sergey ZARITCHNY
--		<sergey.zaritchny@opencascade.com>
---Copyright:	Open CasCade SA 2007

class AsciiStringRetrievalDriver from MDataStd inherits ARDriver from MDF

	---Purpose: Retrieval driver of AsciiString attribute

uses
    RRelocationTable from MDF,
    Attribute        from PDF,
    Attribute        from TDF, 
    MessageDriver    from CDM 
     
is    
    Create(theMessageDriver : MessageDriver from CDM)  -- Version 0
    returns mutable AsciiStringRetrievalDriver from MDataStd;
    

    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type: AsciiString from PDataStd.

    NewEmpty (me)  returns mutable Attribute from TDF;


    Paste(me;
    	  Source     :         Attribute from PDF;
    	  Target     : mutable Attribute from TDF;
    	  RelocTable : RRelocationTable  from MDF);


end AsciiStringRetrievalDriver;
