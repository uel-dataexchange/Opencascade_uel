-- File:	BRepFeat_MakeRevolutionForm.cdl
-- Created:	Tue Oct 14 15:38:43 1997
-- Author:	Olga KOULECHOVA
--		<opt@cleox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


class MakeRevolutionForm from BRepFeat inherits RibSlot from BRepFeat

        ---Purpose: MakeRevolutionForm Generates a surface of
    	-- revolution in the feature as it slides along a
    	-- revolved face in the basis shape.
    	-- The semantics of mechanical features is built
    	-- around giving thickness to a contour. This
    	-- thickness can either be unilateral - on one side
    	-- of the contour - or bilateral - on both sides. As
    	-- in the semantics of form features, the thickness
    	-- is defined by construction of shapes in specific contexts.
    	-- The development contexts differ, however,in
    	-- case of mechanical features. Here they include extrusion:
    	-- -   to a limiting face of the basis shape
    	-- -   to or from a limiting plane
    	-- -   to a height.
        
uses Shape                     from TopoDS,
     Face                      from TopoDS,
     Wire                      from TopoDS,
     Edge                      from TopoDS,
     DataMapOfShapeListOfShape from TopTools,
     Dir                       from gp,
     Ax1                       from gp,
     Vec                       from gp,
     DataMapOfShapeShape       from TopTools,
     ListOfShape               from TopTools,
     SequenceOfCurve           from TColGeom,
     Curve                     from Geom,
     Plane                     from Geom,
     Pnt                       from gp,
     StatusError               from BRepFeat
     
raises ConstructionError from Standard

is


    Create

    	returns MakeRevolutionForm from BRepFeat;
	---Purpose: initializes the linear form class.
	---C++: inline

    Create(Sbase     : Shape   from TopoDS;
	   W         : Wire    from TopoDS;
    	   Plane     : Plane   from Geom; 
	   Axis      : Ax1     from gp;
    	   Height1   : Real    from Standard;
    	   Height2   : Real    from Standard;
    	   Fuse      : Integer from Standard; 
           Sliding   : in out Boolean from Standard)
    
	---Purpose: a contour W, a shape Sbase and a plane P are initialized to serve as
    	--   the basic elements in the construction of the rib or groove. The axis Axis of the
    	--   revolved surface in the basis shape defines the feature's axis of revolution.
    	--   Height1 and Height2 may be used as limits to the construction of the feature.
    	-- Fuse offers a choice between:
    	-- -   removing matter with a Boolean cut using the setting 0 in case of the groove
    	-- -   adding matter with Boolean fusion using the setting 1 in case of the rib.
    		---C++: inline
    	    	returns MakeRevolutionForm from BRepFeat;


    Init(me: in out;  Sbase     : Shape   from TopoDS;
	              W         : Wire    from TopoDS;
	              Plane     : Plane   from Geom; 
	    	      Axis      : Ax1     from gp;
	       	      Height1   : Real    from Standard;	 
	       	      Height2   : Real    from Standard;	 
    	              Fuse      : Integer from Standard; 
                      Sliding   : in out Boolean from Standard)
    
    	is static;
    	---Purpose: Initializes this construction algorithm
    	-- A contour W, a shape Sbase and a plane P are initialized to serve as the basic elements
    	-- in the construction of the rib or groove. The axis Axis of the revolved surface in the basis
    	-- shape defines the feature's axis of revolution. Height1 and Height2 may be
    	-- used as limits to the construction of the feature.
    	-- Fuse offers a choice between:
    	-- -   removing matter with a Boolean cut using the setting 0 in case of the groove
    	-- -   adding matter with Boolean fusion using the setting 1 in case of the rib.
        
    Add(me: in out; E: Edge from TopoDS; OnFace: Face from TopoDS)

	---Purpose: Indicates that the edge <E> will slide on the face
	-- <OnFace>. Raises ConstructionError  if the  face does not belong to the
	-- basis shape, or the edge to the prismed shape.
    	raises ConstructionError from Standard
	
	is static;



    Perform(me: in out)
    
    	is static;
    	---Purpose: Performs a prism from the wire to the plane
    	-- along the basis shape S. Reconstructs the feature topologically.


    Propagate(me: in out; L: in out ListOfShape from TopTools;
    	    	    	  F: Face from TopoDS;
    	    	    	  FPoint, LPoint:   Pnt from gp; 
    	    	    	  falseside : in out Boolean from Standard)
	returns Boolean from Standard
	is static;


fields

    myAxe      : Ax1                       from gp;
    myHeight1  : Real                      from Standard;
    myHeight2  : Real                      from Standard;
    mySliding  : Boolean                   from Standard;
    myPln      : Plane                     from Geom;    
    myBnd      : Real                      from Standard;
    mySlface   : DataMapOfShapeListOfShape from TopTools;
    myListOfEdges : ListOfShape            from TopTools;
    myTol      : Real                      from Standard;
    myAngle1   : Real                      from Standard;
    myAngle2   : Real                      from Standard;

end MakeRevolutionForm;



