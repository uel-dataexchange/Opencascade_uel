-- File:	MDataStd_TreeNodeRetrievalDriver.cdl
-- Created:	Thu Jun 17 12:10:22 1999
-- Author:	Vladislav ROMASHKO
--		<vro@flox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999

class TreeNodeRetrievalDriver from MDataStd inherits ARDriver from MDF


uses 
     
     RRelocationTable from MDF,
     Attribute        from PDF,
     Attribute        from TDF, 
     MessageDriver    from CDM

is
 
    Create (theMessageDriver : MessageDriver from CDM) 
     returns mutable TreeNodeRetrievalDriver from MDataStd;
    
    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;

    NewEmpty (me)  returns mutable Attribute from TDF;

    Paste(me;
    	  Source     :         Attribute from PDF;
    	  Target     : mutable Attribute from TDF;
    	  RelocTable : RRelocationTable  from MDF);

end TreeNodeRetrievalDriver;
