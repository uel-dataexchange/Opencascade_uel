-- File:        ApprovalStatus.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWApprovalStatus from RWStepBasic

	---Purpose : Read & Write Module for ApprovalStatus

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ApprovalStatus from StepBasic

is

	Create returns RWApprovalStatus;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ApprovalStatus from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : ApprovalStatus from StepBasic);

end RWApprovalStatus;
