--
-- File      :  RightAngularWedge.cdl
-- Created   :  Sat 9 Jan 1993
-- Author    : CKY / Contract Toubro-Larsen ( SIVA )
--
---Copyright : MATRA-DATAVISION  1993
--

class RightAngularWedge from IGESSolid  inherits IGESEntity


        ---Purpose: defines RightAngularWedge, Type <152> Form Number <0>
        --          in package IGESSolid
        --          A right angular wedge is a triangular/trapezoidal prism

uses

        Pnt             from gp,
        Dir             from gp,
        XYZ             from gp

is

        Create returns mutable RightAngularWedge;

        Init (me         : mutable;
              aSize      : XYZ;
              lowX       : Real;
              aCorner    : XYZ;
              anXAxis    : XYZ;
              anZAxis    : XYZ);
        ---Purpose : This method is used to set the fields of the class
        --           RightAngularWedge
        --       - aSize    : the lengths along the local axes
        --       - lowX     : the length at the smaller X-side
        --       - aCorner  : the corner point coordinates
        --                    default (0,0,0)
        --       - anXAxis  : the unit vector defining local X-axis
        --                    default (1,0,0)
        --       - anZAxis  : the unit vector defining local Z-axis
        --                    default (0,0,1)
    
        Size(me) returns XYZ;
        ---Purpose : returns the size

        XBigLength (me) returns Real;
        ---Purpose : returns the length along the local X-axis

        XSmallLength (me) returns Real;
        ---Purpose : returns the smaller length along the local X-direction at Y=LY

        YLength (me) returns Real;
        ---Purpose : returns the length along the local Y-axis

        ZLength (me) returns Real;
        ---Purpose : returns the length along the local Z-axis

        Corner (me) returns Pnt;
        ---Purpose : returns the corner point coordinates

        TransformedCorner (me) returns Pnt;
        ---Purpose : returns the corner point coordinates after applying
        -- TransformationMatrix

        XAxis (me) returns Dir;
        ---Purpose : returns the direction defining the local X-axis

        TransformedXAxis (me) returns Dir;
        ---Purpose : returns the direction defining the local X-axis
        -- after applying the TransformationMatrix

        YAxis (me) returns Dir;
        ---Purpose : returns the direction defining the local Y-axis
        -- it is got by taking the cross product of ZAxis and XAxis

        TransformedYAxis (me) returns Dir;
        ---Purpose : returns the direction defining the local Y-axis
        -- after applying the TransformationMatrix

        ZAxis (me) returns Dir;
        ---Purpose : returns the direction defining the local Z-axis

        TransformedZAxis (me) returns Dir;
        ---Purpose : returns the direction defining the local Z-axis
        -- after applying the TransformationMatrix

fields

--
-- Class    : IGESSolid_RightAngularWedge
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class RightAngularWedge.
--
-- Reminder : A RightAngularWedge instance is defined by :
--            a vertex at (X1,Y1,Z1) and three orthogonal edges lying
--            along the local +X, +Y and +Z axes. The local X and Z axes
--            are defined by a unit vector along the axes.

        theSize          : XYZ;     
            -- the lengths along the local axes

        theXSmallLength  : Real;
            -- the length of X-direction at Y = LY

        theCorner        : XYZ;
            -- the corner point coordinates

        theXAxis         : XYZ;
            -- the unit vector along the local X-direction

        theZAxis         : XYZ;
            -- the unit vector along the local Z-direction

end RightAngularWedge;
