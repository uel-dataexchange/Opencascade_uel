-- File:        Polyline.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPolyline from RWStepGeom

	---Purpose : Read & Write Module for Polyline

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Polyline from StepGeom,
     EntityIterator from Interface

is

	Create returns RWPolyline;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Polyline from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : Polyline from StepGeom);

	Share(me; ent : Polyline from StepGeom; iter : in out EntityIterator);

end RWPolyline;
