-- File:	RWStepRepr_RWConfigurationEffectivity.cdl
-- Created:	Fri Nov 26 16:26:36 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWConfigurationEffectivity from RWStepRepr

    ---Purpose: Read & Write tool for ConfigurationEffectivity

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ConfigurationEffectivity from StepRepr

is
    Create returns RWConfigurationEffectivity from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ConfigurationEffectivity from StepRepr);
	---Purpose: Reads ConfigurationEffectivity

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ConfigurationEffectivity from StepRepr);
	---Purpose: Writes ConfigurationEffectivity

    Share (me; ent : ConfigurationEffectivity from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWConfigurationEffectivity;
