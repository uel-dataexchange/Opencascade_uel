-- File:	StepData_StepDumper.cdl
-- Created:	Mon Mar 14 10:38:08 1994
-- Author:	Christian CAILLET
--		<cky@ecolox>
---Copyright:	 Matra Datavision 1994


class StepDumper  from StepData

    ---Purpose : Provides a way to dump entities processed through STEP, with
    --           these features :
    --           - same form as for writing a STEP File (because it is clear
    --             and compact enough, even if the names of the fields do not
    --             appear) : thus, no additionnal resource is required
    --           - possibility to look for an entity itself (only its Type or
    --             with its content), an entity and it shared items (one level)
    --             or all the entities its refers to, directly or recursively.

uses Messenger from Message, Transient, Protocol from StepData, StepModel,
     GeneralLib, StepWriter, WriterLib

raises InterfaceMismatch

is

    Create (amodel : StepModel; protocol : Protocol from StepData; mode : Integer = 0)
    	    returns StepDumper;
    ---Purpose : Creates a StepDumper, able to work on a given StepModel
    --           (which defines the total scope for dumping entities) and
    --           a given Protocol from Step (which defines the authorized
    --           types to be dumped)
    --           <mode> commands what is to be displayed (number or label)
    --           0 for number (and corresponding labels  are displayed apart)
    --           1 for label  (and corresponding numbers are displayed apart)
    --           2 for label without anymore

    StepWriter (me : in out) returns StepWriter  is static;
    ---Purpose : Gives an access to the tool which is used to work : this allow
    --           to acts on some parameters : Floating Format, Scopes ...
    ---C++ : return &

    Dump (me : in out; S : Messenger from Message; ent : Transient; level : Integer)
        returns Boolean
    ---Purpose : Dumps a Entity on an Messenger. Returns True if
    --           sucess, False, if the entity to dump has not been recognized
    --           by the Protocol. <level> can have one of these values :
    --           - 0 : prints the TYPE only, as known in STEP Files (StepType)
    --             If <ent> has not been regognized by the Protocol, or if its
    --             type is Complex, the StepType is replaced by the display of
    --             the cdl type. Complex Type are well processed by level 1.
    --           - 1 : dumps the entity, completely (whatever it has simple or
    --             complex type) but alone.
    --           - 2 : dumps the entity completely, plus the item its refers to
    --                 at first level (a header message designates the starting
    --                 entity of the dump) <Lists Shared and Implied>
    --           - 3 : dumps the entity and its refered items at any levels
    --           
    --           For levels 1,2,3, the numbers displayed (form #nnn) are the
    --           numbers of the corresponding entities in the Model
    	raises InterfaceMismatch;
    --           Errors come from StepWriter, they especially occur when an
    --           entity does not come from the starting Model.
    --           Level 0 accepts an entity which does not come from the Model.

    Dump (me : in out; S : Messenger from Message; num : Integer; level : Integer)
        returns Boolean
    ---Purpose : Works as Dump with a Transient, but directly takes the
    --           entity designated by its number in the Model
    --           Returns False, also if <num> is out of range
    	raises InterfaceMismatch;
    --           Errors : same as above

fields

    themodel  : StepModel;
    theslib   : GeneralLib;
    thewlib   : WriterLib;
    thewriter : StepWriter;

end StepDumper;
