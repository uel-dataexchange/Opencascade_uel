-- File:	RWStepRepr_RWDerivedShapeAspect.cdl
-- Created:	Wed Jun  4 14:17:23 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWDerivedShapeAspect from RWStepRepr

    ---Purpose: Read & Write tool for DerivedShapeAspect

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    DerivedShapeAspect from StepRepr

is
    Create returns RWDerivedShapeAspect from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : DerivedShapeAspect from StepRepr);
	---Purpose: Reads DerivedShapeAspect

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: DerivedShapeAspect from StepRepr);
	---Purpose: Writes DerivedShapeAspect

    Share (me; ent : DerivedShapeAspect from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWDerivedShapeAspect;
