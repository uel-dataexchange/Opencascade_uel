-- File:	RWStepAP214_RWAppliedOrganizationAssignment.cdl
-- Created:	Fri Mar 12 12:03:16 1999
-- Author:	data exchange team
--		<det@androx.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class RWAppliedOrganizationAssignment from RWStepAP214 

	---Purpose: Read & Write Module for AppliedOrganizationAssignment

uses
     Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     AppliedOrganizationAssignment from StepAP214,
     EntityIterator from Interface

is
    	Create returns RWAppliedOrganizationAssignment;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable AppliedOrganizationAssignment from StepAP214);

	WriteStep (me; SW : in out StepWriter; ent : AppliedOrganizationAssignment from StepAP214);

	Share(me; ent : AppliedOrganizationAssignment from StepAP214; iter : in out EntityIterator);

end RWAppliedOrganizationAssignment;
