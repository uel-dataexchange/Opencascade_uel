-- File     : Prs2d_Angle.cdl
-- Created  : February  2000
-- Author   : Tanya COOL
---Copyright: Matra Datavision 2000

class Angle from Prs2d inherits Dimension from Prs2d

 ---Purpose: Constructs the primitive Angle

uses

	Drawer		   from Graphic2d,
	GraphicObject	   from Graphic2d,
	Pnt2d              from gp,
	Length             from Quantity,
	ExtendedString     from TCollection,
	ArrowSide          from Prs2d,
	TypeOfArrow        from Prs2d,
        FStream            from Aspect 

raises

	CircleDefinitionError	from Graphic2d

is
	Create( aGraphicObject: GraphicObject  from Graphic2d;
	        anAttachPnt1  : Pnt2d          from gp;
		anAttachPnt2  : Pnt2d          from gp;
            	anAttachPnt3  : Pnt2d          from gp;
            	aRadius       : Length         from Quantity;
	        aText         : ExtendedString from TCollection;
	        aTxtScale     : Real           from Standard = 3.0;
	        anArrAngle    : Real           from Standard = 15.0;
	        anArrLength   : Real           from Standard = 10.0;
	        anArrType     : TypeOfArrow    from Prs2d = Prs2d_TOA_OPENED;
	        anArrow       : ArrowSide      from Prs2d = Prs2d_AS_BOTHAR;
	        IsReverseArrow: Boolean        from Standard = Standard_False )

	returns mutable Angle from Prs2d;

	---Purpose: create an angle:
    	--          between the line defined by the points
    	--          anAttachtPnt1 and anAttachPnt2 and
    	--          the line defined by the points
    	--          anAttachPnt1 and anAttachPnt3
    	--          Radius of this angle is the distance 
    	--          between <anAttachPnt1> and <anOffsetPoint> points.
    	--          <anArrAngle> in degree
   
        --------------------------------------
	-- Category: Inquire methods
	--------------------------------------
    
    Values( me; aPnt1, aPnt2, aPnt3: out Pnt2d from gp; 
            aRad: out Length from Quantity ); 
    	---Level: Internal
    	---Purpose: allows to get the properties of the angle
    
    CalcTxtPos(me:mutable; theFromAbs: Boolean 
    	        from Standard=Standard_False) 
	---C++: inline
	is redefined protected;
    
	--------------------------------------
	-- Category: Draw and Pick
	--------------------------------------

    Draw( me : mutable; aDrawer: Drawer from Graphic2d )
	is static protected;
	---Level: Internal
	---Purpose: Draws the angle <me>.

    DrawElement( me : mutable; aDrawer: Drawer from Graphic2d;
                 anIndex: Integer from Standard)
        is redefined protected;
    	---Level: Internal
    	---Purpose: Draws element <anIndex> of the angle <me>.

    DrawVertex( me : mutable; aDrawer: Drawer from Graphic2d;
                anIndex: Integer from Standard)
        is redefined protected;
    	---Level: Internal
    	---Purpose: Draws vertex <anIndex> of the angle <me>.

    Pick( me : mutable; X, Y: ShortReal from Standard;
	  aPrecision: ShortReal from Standard;
	  aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard
	is static protected;
	---Level: Internal
	---Purpose: Returns Standard_True if the angle <me> is picked,
	--	    Standard_False if not.

    Save( me; aFStream: in out FStream from Aspect ) is virtual;
														
fields
 
	myCentX          : ShortReal         from Standard;
	myCentY          : ShortReal         from Standard;
	myRad            : ShortReal         from Standard;
        myFAngle         : ShortReal         from Standard;
    	mySAngle         : ShortReal         from Standard;
	
end Angle from Prs2d;
