-- File:	IGESGeom_ToolOffsetCurve.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolOffsetCurve  from IGESGeom

    ---Purpose : Tool to work on a OffsetCurve. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses OffsetCurve from IGESGeom,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolOffsetCurve;
    ---Purpose : Returns a ToolOffsetCurve, ready to work


    ReadOwnParams (me; ent : mutable OffsetCurve;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : OffsetCurve;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : OffsetCurve;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a OffsetCurve <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable OffsetCurve) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a OffsetCurve
    --           (if OffsetType is not 3, OffsetFunction is cleared)

    DirChecker (me; ent : OffsetCurve) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : OffsetCurve;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : OffsetCurve; entto : mutable OffsetCurve;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : OffsetCurve;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolOffsetCurve;
