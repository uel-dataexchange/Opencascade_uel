---Copyright:	 Matra Datavision 1992
---Version: 

---History:
--  Version	Date         Purpose
--              18/12/92     Creation   

generic class HIndexedDataMap from PCollection ( Key      as Storable;
		            	            Item     as Storable;
			    	    	    KeyHash  as Hash(Key)
    	    	    	    	    	 )
	    
---Purpose: The HIndexedDataMap is a hashed set of objects of Type Key, called 
-- Keys. Keys can be inserted in the Map but not removed. The Map 
-- keeps the number of keys called NbKeys. Each time a Key is
-- inserted the Map tests if this Key is already in the Map. If 
-- it is, nothing is done. If not, NbKeys is incremented and it's 
-- value is bound to the Key and called the Index.
-- 
-- The Map provides methods to inquire the Index of a Key and to 
-- retrieve a Key from an Index in the range 1..NbKeys.
-- 
-- Another Datum of the type Item can be stored with the Key. The 
-- Item can be retrieved from the Key and from the Index of the
-- Key. The Item stored with a Key can be modified.

inherits Persistent from Standard

raises

    OutOfRange from Standard
    

class IndexedDataMapNode from PCollection inherits PManaged from PMMgt

---Purpose: This class is used in the implementation of the IndexedDataMap class. 
-- It stores three elements : a Key, an Item and an Integer Index. 
-- It  also stores two references to IndexedDataMapNode objects, 
-- IndexedDataMapNode are used to make lists in the Hashed IndexedDataMap.

is

    Create(aKey : Key; Index : Integer; anItem : Item; NextKey,NextIndex
    	: IndexedDataMapNode )returns mutable IndexedDataMapNode;
    ---Purpose: Creates a IndexedDataMapNode;

    Set(me : mutable; aKey : Key; Index : Integer; anItem : Item; 
    	    NextK,NextI : IndexedDataMapNode) is static;
    ---Level: Internal
    ---Purpose: Sets the values of <me>.

    SetItem ( me : mutable; anItem : Item) is static;
    ---Level: Internal
    ---Purpose: Sets the item.
    
    SetNextKey ( me : mutable ; aNode : IndexedDataMapNode ) is static;
    ---Level: Internal
    ---Purpose: Sets the next node of Key hashed list.

    SetNextIndex ( me : mutable ; aNode : IndexedDataMapNode ) is static;
    ---Level: Internal
    ---Purpose: Sets the next node of Key hashed list.

    GetKey ( me ) returns any Key is static;
    ---Level: Internal
    ---Purpose: Returns the key.
    
    Index ( me ) returns Integer is static;
    ---Level: Internal
    ---Purpose: Returns the index.
    
    GetItem ( me ) returns any Item is static;
    ---Level: Internal
    ---Purpose: Returns the item.
    
    IndexAndItem(me; Index : out Integer; theItem : out any Item) is static;
    ---Level: Internal
    ---Purpose: Returns index and item.
    
    KeyAndItem(me; theKey : out any Key; theItem : out any Item) is static;
    ---Level: Internal
    ---Purpose: Returns key and item.
    
    NextKey ( me ) returns any IndexedDataMapNode is static;
    ---Level: Internal
    ---Purpose: Returns the next node of Key hashed list.

    NextIndex ( me ) returns any IndexedDataMapNode is static;
    ---Level: Internal
    ---Purpose: Returns the next node of Index hashed list.

fields

    myKey       : Key;
    myIndex     : Integer;
    myItem      : Item;
    myNextKey   : IndexedDataMapNode;
    myNextIndex : IndexedDataMapNode;

end IndexedDataMapNode;
    
class ArrayIndexedDataMap instantiates 
                       HArray1 from PCollection (IndexedDataMapNode);
    
is

    Create ( NbBuckets : Integer; fhKey : KeyHash ) returns mutable HIndexedDataMap;
    ---Purpose: Creates an empty HIndexedDataMap, NbBuckets is an estimation of the
    -- number of Keys that will be stored in the Map. It is not 
    -- limited, but a too small number may reduce performance.

    NbBuckets ( me ) returns Integer;
    ---Level: Public
    ---Purpose: Returns the number of entries in the indexed map.

    NbKeys(me) returns Integer;
    ---Level: Public
    ---Purpose: Returns the number of Keys stored in the Map.
    
    Bind(me : mutable ; aKey : Key; anItem : Item; OverWrite : Boolean ) 
    	returns Integer;
    ---Level: Public
    ---Purpose: Adds a new Key and returns the Index. 
    -- If the Key is new in the Map the Item is bound with the Key. 
    -- If the Key is already present the Item replaces the existing
    -- Item if Overwrite is True.
    
    FindIndex ( me ; aKey : Key ) returns Integer;
    ---Level: Public
    ---Purpose: Returns the Index of the Key in the Map. If the Key is not 
    -- stored the returned Index is 0.
    
    FindKey ( me ; Index : Integer ) returns any Key
    ---Level: Public
    ---Purpose: Returns the Key stored with the Index, Index must be in the 
    -- range 1..NbKeys.
    raises OutOfRange from Standard;
    
    FindItemFromKey ( me ; aKey : Key ) returns any Item
    ---Level: Public
    ---Purpose: Returns the Item stored with the Key <aKey>.
    ---Trigger: An exception is raised if the key <aKey> is not stored in the Map.
    raises OutOfRange from Standard;
    
    FindItemFromIndex ( me ; Index : Integer ) returns any Item
    ---Level: Public
    ---Purpose: Returns the Item stored with the index <Index>. This  is 
    -- similar to but faster than K = GetKey(Index); GetItem(K,I)
    ---Trigger: An exception is raised if <Index> is not in the range 1..NbKeys.
    raises OutOfRange from Standard;
    
    FindIndexAndItem(me; aKey : Key; Index : out Integer; theItem : out Item)
    ---Level: Public
    ---Purpose: Returns the index and the item stored with the Key <aKey>.
    ---Trigger: An exception is raised if the key <aKey> is not stored in the Map.
    raises OutOfRange from Standard;
    
    FindKeyAndItem(me; Index : Integer; theKey : out Key; theItem : out Item)
    ---Level: Public
    ---Purpose: Returns the key and the item stored with the index <Index>.
    ---Trigger: An exception is raised if <Index> is not in the range 1..NbKeys.
    raises OutOfRange from Standard;
    
    SetItemToKey(me : mutable; aKey : Key; anItem : Item)
    ---Level: Public
    ---Purpose: Modifies the item stored with the key <aKey>.
    ---Trigger: An exception is raised if the key <aKey> is not stored in the Map.
    raises OutOfRange from Standard;
    
    SetItemToIndex(me : mutable; Index : Integer; anItem : Item)
    ---Level: Public
    ---Purpose: Modifies the item stored with the index <Index>.
    ---Trigger: An exception is raised if <Index> is not in the range 1..NbKeys.
    raises OutOfRange from Standard;

    Clear ( me : mutable );
    ---Level: Public
    ---Purpose: Clears the Map content.
    
    IsBound ( me ; aKey : Key) returns Boolean;
    ---Level: Public
    ---Purpose: Returns True if an element is bound by <aKey>.
    
    LocateKey(me; aKey : Key) returns any IndexedDataMapNode
    ---Level: Internal
    ---Purpose: Returns the node containing <aKey>.
    is static private;
    
    LocateIndex(me; Index : Integer) returns any IndexedDataMapNode
    ---Level: Internal
    ---Purpose: Returns the node containing <Index>.
    is static private;
    
fields

    myNumber       : Integer;
    myKeyHash      : KeyHash;
    myArrayKey     : ArrayIndexedDataMap;
    myArrayIndices : ArrayIndexedDataMap;
    
end HIndexedDataMap;




