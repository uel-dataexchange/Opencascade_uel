-- File:        ContextDependentOverRidingStyledItem.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWContextDependentOverRidingStyledItem from RWStepVisual

	---Purpose : Read & Write Module for ContextDependentOverRidingStyledItem

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ContextDependentOverRidingStyledItem from StepVisual,
     EntityIterator from Interface

is

	Create returns RWContextDependentOverRidingStyledItem;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ContextDependentOverRidingStyledItem from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : ContextDependentOverRidingStyledItem from StepVisual);

	Share(me; ent : ContextDependentOverRidingStyledItem from StepVisual; iter : in out EntityIterator);

end RWContextDependentOverRidingStyledItem;
