-- File:        SiUnitAndPlaneAngleUnit.cdl
-- Created:     Mon Dec  4 12:02:36 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSiUnitAndPlaneAngleUnit from RWStepBasic

	---Purpose : Read & Write Module for SiUnitAndPlaneAngleUnit

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SiUnitAndPlaneAngleUnit from StepBasic

is

    Create returns RWSiUnitAndPlaneAngleUnit;

    ReadStep (me; data : StepReaderData; num : Integer;
	      ach : in out Check; ent : mutable SiUnitAndPlaneAngleUnit from StepBasic);

    WriteStep (me; SW : in out StepWriter; ent : SiUnitAndPlaneAngleUnit from StepBasic);

	  
end RWSiUnitAndPlaneAngleUnit;
