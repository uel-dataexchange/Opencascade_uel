-- File:        OrdinalDate.cdl
-- Created:     Fri Dec  1 11:11:22 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class OrdinalDate from StepBasic 

inherits Date from StepBasic 

uses

	Integer from Standard
is

	Create returns mutable OrdinalDate;
	---Purpose: Returns a OrdinalDate


	Init (me : mutable;
	      aYearComponent : Integer from Standard) is redefined;

	Init (me : mutable;
	      aYearComponent : Integer from Standard;
	      aDayComponent : Integer from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetDayComponent(me : mutable; aDayComponent : Integer);
	DayComponent (me) returns Integer;

fields

	dayComponent : Integer from Standard;

end OrdinalDate;
