-- File:	RWStepShape_RWShapeDimensionRepresentation.cdl
-- Created:	Tue Apr 18 16:42:59 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWShapeDimensionRepresentation from RWStepShape

    ---Purpose: Read & Write tool for ShapeDimensionRepresentation

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ShapeDimensionRepresentation from StepShape

is
    Create returns RWShapeDimensionRepresentation from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ShapeDimensionRepresentation from StepShape);
	---Purpose: Reads ShapeDimensionRepresentation

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ShapeDimensionRepresentation from StepShape);
	---Purpose: Writes ShapeDimensionRepresentation

    Share (me; ent : ShapeDimensionRepresentation from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWShapeDimensionRepresentation;
