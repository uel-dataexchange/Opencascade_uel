-- File:	GeomToIGES_GeomPoint.cdl
-- Created:	Wed Nov 16 14:24:57 1994
-- Author:	Marie Jose MARTZ
--		<mjm@minox>
---Copyright:	 Matra Datavision 1994

class GeomPoint from GeomToIGES inherits GeomEntity from GeomToIGES

    ---Purpose: This class implements the transfer of the Point Entity from Geom
    --          to IGES . These are :
    --          . Point
    --              * CartesianPoint 

  
uses

    Point          from Geom,
    CartesianPoint from Geom,
    Point          from IGESGeom,
    GeomEntity     from GeomToIGES
     
is 
    
    Create returns GeomPoint from GeomToIGES;


    Create(GE : GeomEntity from GeomToIGES)  
    	 returns GeomPoint from GeomToIGES;
    ---Purpose : Creates a tool GeomPoint ready to run and sets its
    --         fields as GE's.

    TransferPoint            (me    : in out;
                              start : Point from Geom)
    	 returns mutable Point from IGESGeom;
    ---Purpose :  Transfert  a  Point from Geom to IGES. If this
    --            Entity could not be converted, this member returns a NullEntity.

    TransferPoint            (me    : in out;
                              start : CartesianPoint from Geom)
    	 returns mutable Point from IGESGeom;
    ---Purpose :  Transfert  a  CartesianPoint from Geom to IGES. If this
    --            Entity could not be converted, this member returns a NullEntity.


end GeomPoint;


