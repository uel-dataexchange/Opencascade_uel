-- File:        RepresentationItem.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWRepresentationItem from RWStepRepr

	---Purpose : Read & Write Module for RepresentationItem

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     RepresentationItem from StepRepr

is

	Create returns RWRepresentationItem;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable RepresentationItem from StepRepr);

	WriteStep (me; SW : in out StepWriter; ent : RepresentationItem from StepRepr);

end RWRepresentationItem;
