-- File:	IGESGeom_ToolTrimmedSurface.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolTrimmedSurface  from IGESGeom

    ---Purpose : Tool to work on a TrimmedSurface. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses TrimmedSurface from IGESGeom,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolTrimmedSurface;
    ---Purpose : Returns a ToolTrimmedSurface, ready to work


    ReadOwnParams (me; ent : mutable TrimmedSurface;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : TrimmedSurface;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : TrimmedSurface;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a TrimmedSurface <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : TrimmedSurface) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : TrimmedSurface;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : TrimmedSurface; entto : mutable TrimmedSurface;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : TrimmedSurface;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolTrimmedSurface;
