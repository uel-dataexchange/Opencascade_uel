--
-- File      :  SelectedComponent.cdl
-- Created   :  Sat 9 Jan 1993
-- Author    : CKY / Contract Toubro-Larsen ( SIVA )
--
---Copyright : MATRA-DATAVISION  1993
--

class SelectedComponent from IGESSolid  inherits IGESEntity

        ---Purpose: defines SelectedComponent, Type <182> Form Number <0>
        --          in package IGESSolid
        --          The Selected Component entity provides a means of
        --          selecting one component of a disjoint CSG solid

uses

        BooleanTree     from IGESSolid,
        XYZ             from gp,
        Pnt             from gp

is

        Create returns mutable SelectedComponent;

        -- Specific Methods pertaining to the class

        Init (me        : mutable;
              anEntity  : BooleanTree;
              selectPnt : XYZ);
        ---Purpose : This method is used to set the fields of the class
        --           SelectedComponent
        --       - anEntity  : the Boolean tree entity
        --       - selectPnt : Point in or on the desired component

        Component(me) returns BooleanTree;
        ---Purpose : returns the Boolean tree entity

        SelectPoint(me) returns Pnt;
        ---Purpose : returns the point on/in the selected component

        TransformedSelectPoint(me) returns Pnt;
        ---Purpose : returns the point on/in the selected component
        -- after applying TransformationMatrix

fields

--
-- Class    : IGESSolid_SelectedComponent
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class SelectedComponent.
--
-- Reminder : A SelectedComponent instance is defined by :
--            a pointer to the Boolean Tree entity(Entity) and the X, Y
--            and Z components (X,Y,Z) of a selected point.

        theEntity      : BooleanTree;
            -- the desired boolean tree entity

        theSelectPoint : XYZ;
            -- the X, Y and Z coordinates of the point

end SelectedComponent;
