-- File:        Loop.cdl
-- Created:     Mon Dec  4 12:02:27 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWLoop from RWStepShape

	---Purpose : Read & Write Module for Loop

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Loop from StepShape

is

	Create returns RWLoop;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Loop from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : Loop from StepShape);

end RWLoop;
