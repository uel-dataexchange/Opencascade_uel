-- File:	StepToGeom_MakeCurve.cdl
-- Created:	Mon Jun 21 10:14:42 1993
-- Author:	Martine LANGLOIS
---Copyright:	 Matra Datavision 1993

class MakeCurve from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          class Curve from StepGeom which
    --          describes a Curve from prostep and Curve from Geom. 
    --          As Curve is an abstract class
    --          this class an access to the sub-class required.

uses Curve from Geom,
     Curve from StepGeom

is 

    Convert ( myclass; SC : Curve from StepGeom;
                       CC : out Curve from Geom )
    returns Boolean from Standard;

end MakeCurve;
