-- File:        PresentationSizeAssignmentSelect.cdl
-- Created:     Fri Dec  1 11:11:11 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class PresentationSizeAssignmentSelect from StepVisual inherits SelectType from StepData

	-- <PresentationSizeAssignmentSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : PresentationView, PresentationArea, AreaInSet

uses

	PresentationView,
	PresentationArea,
	AreaInSet
is

	Create returns PresentationSizeAssignmentSelect;
	---Purpose : Returns a PresentationSizeAssignmentSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a PresentationSizeAssignmentSelect Kind Entity that is :
	--        1 -> PresentationView
	--        2 -> PresentationArea
	--        3 -> AreaInSet
	--        0 else

	PresentationView (me) returns any PresentationView;
	---Purpose : returns Value as a PresentationView (Null if another type)

	PresentationArea (me) returns any PresentationArea;
	---Purpose : returns Value as a PresentationArea (Null if another type)

	AreaInSet (me) returns any AreaInSet;
	---Purpose : returns Value as a AreaInSet (Null if another type)


end PresentationSizeAssignmentSelect;

