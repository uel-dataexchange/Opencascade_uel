-- File:	StepDimTol_GeometricToleranceRelationship.cdl
-- Created:	Wed Jun  4 13:34:35 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class GeometricToleranceRelationship from StepDimTol
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity GeometricToleranceRelationship

uses
    HAsciiString from TCollection,
    GeometricTolerance from StepDimTol

is
    Create returns GeometricToleranceRelationship from StepDimTol;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       aDescription: HAsciiString from TCollection;
                       aRelatingGeometricTolerance: GeometricTolerance from StepDimTol;
                       aRelatedGeometricTolerance: GeometricTolerance from StepDimTol);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

    RelatingGeometricTolerance (me) returns GeometricTolerance from StepDimTol;
	---Purpose: Returns field RelatingGeometricTolerance
    SetRelatingGeometricTolerance (me: mutable; RelatingGeometricTolerance: GeometricTolerance from StepDimTol);
	---Purpose: Set field RelatingGeometricTolerance

    RelatedGeometricTolerance (me) returns GeometricTolerance from StepDimTol;
	---Purpose: Returns field RelatedGeometricTolerance
    SetRelatedGeometricTolerance (me: mutable; RelatedGeometricTolerance: GeometricTolerance from StepDimTol);
	---Purpose: Set field RelatedGeometricTolerance

fields
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection;
    theRelatingGeometricTolerance: GeometricTolerance from StepDimTol;
    theRelatedGeometricTolerance: GeometricTolerance from StepDimTol;

end GeometricToleranceRelationship;
