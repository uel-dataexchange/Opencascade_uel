-- File:	MXCAFDoc_DimTolRetrievalDriver.cdl
-- Created:	Wed Dec 10 09:48:30 2008
-- Author:	Pavel TELKOV
--		<ptv@valenox>
---Copyright:	 Open CASCADE 2008

class DimTolRetrievalDriver from MXCAFDoc inherits ARDriver from MDF

	---Purpose: 
uses
    RRelocationTable from MDF,
    Attribute        from PDF,
    Attribute        from TDF,
    MessageDriver    from CDM

is
    Create (theMsgDriver : MessageDriver from CDM)
    returns mutable DimTolRetrievalDriver from MXCAFDoc;
	---Purpose: Returns mutable DimTolRetrievalDriver from MXCAFDoc;

    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
    ---Purpose: Returns the type: XCAFDoc_DimTol

    NewEmpty (me)  returns mutable Attribute from TDF;

    Paste(me;
    	  Source     :         Attribute from PDF;
    	  Target     : mutable Attribute from TDF;
    	  RelocTable : RRelocationTable from MDF);

end DimTolRetrievalDriver from MXCAFDoc;
