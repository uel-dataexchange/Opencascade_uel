-- File:	RWStepBasic_RWActionMethod.cdl
-- Created:	Fri Nov 26 16:26:29 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWActionMethod from RWStepBasic

    ---Purpose: Read & Write tool for ActionMethod

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ActionMethod from StepBasic

is
    Create returns RWActionMethod from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ActionMethod from StepBasic);
	---Purpose: Reads ActionMethod

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ActionMethod from StepBasic);
	---Purpose: Writes ActionMethod

    Share (me; ent : ActionMethod from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWActionMethod;
