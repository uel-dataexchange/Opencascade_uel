-- File:	Geom2d_BoundedCurve.cdl
-- Created:	Wed Mar 24 17:54:32 1993
-- Author:	JCV
--		<fid@sdsun2>
-- Copyright:	 Matra Datavision 1993

---Copyright:   Matra Datavision 1991



deferred class BoundedCurve from Geom2d inherits Curve from Geom2d 

    	--- Purpose : The abstract class BoundedCurve describes the
    	-- common behavior of bounded curves in 2D space. A
    	-- bounded curve is limited by two finite values of the
    	-- parameter, termed respectively "first parameter" and
    	-- "last parameter". The "first parameter" gives the "start
    	-- point" of the bounded curve, and the "last parameter"
    	-- gives the "end point" of the bounded curve.
    	-- The length of a bounded curve is finite.
    	-- The Geom2d package provides three concrete
    	-- classes of bounded curves:
    	-- - two frequently used mathematical formulations of complex curves:
    	--   - Geom2d_BezierCurve,
    	--   - Geom2d_BSplineCurve, and
    	-- - Geom2d_TrimmedCurve to trim a curve, i.e. to
    	--   only take part of the curve limited by two values of
    	--   the parameter of the basis curve.

uses Pnt2d from gp


is

  EndPoint (me)   returns Pnt2d  is deferred;
        --- Purpose : 
        --  Returns the end point of the curve.
        --  The end point is the value of the curve for the 
        --  "LastParameter" of the curve.


  StartPoint (me)  returns Pnt2d   is deferred;
        --- Purpose : 
        --  Returns the start point of the curve.
        --  The start point is the value of the curve for the 
        --  "FirstParameter" of the curve.


end;
