-- File:        PointStyle.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPointStyle from RWStepVisual

	---Purpose : Read & Write Module for PointStyle

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PointStyle from StepVisual,
     EntityIterator from Interface

is

	Create returns RWPointStyle;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PointStyle from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : PointStyle from StepVisual);

	Share(me; ent : PointStyle from StepVisual; iter : in out EntityIterator);

end RWPointStyle;
