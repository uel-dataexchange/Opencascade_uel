-- File:       PlotMgt_PlotterDriver.cdl
-- Created:    25-NOV-98
-- Author:     DCB
---Copyright:  Matra Datavision 1998
-- Updated:	GG 03/10/00 BUC60766 The Close() method can be used for freeing
--		the opened file and must be declared accessible by any client.

deferred class PlotterDriver from PlotMgt inherits Driver from Aspect

uses
  PlaneAngle        from Quantity,
  Factor            from Quantity,
  Ratio             from Quantity,
  Length            from Quantity,
  ColorMap          from Aspect, 
  TypeMap           from Aspect,
  WidthMap          from Aspect, 
  MarkMap           from Aspect, 
  FontMap           from Aspect, 
  ExtendedString    from TCollection,     
  TypeOfText        from Aspect,
  TypeOfColorSpace  from Aspect,
  TypeOfPrimitive   from Aspect,
  PlotMode          from Aspect,
  FStream           from Aspect,
  Plotter           from PlotMgt,
  HListOfMFTFonts   from PlotMgt,
  HArray1OfShortReal from TShort,
  TextManager       from PlotMgt,
  AsciiString       from TCollection,
  Array1OfShortReal from TShort


is
  Initialize (aPlotter    : Plotter from PlotMgt;
      aFileName   : CString from Standard;
      fCreateFile : Boolean from Standard = Standard_False);
      ---Level: Private

  Initialize (aFileName   : CString from Standard;              
      fCreateFile : Boolean from Standard = Standard_False);
      ---Level: Private

  BeginDraw (me: mutable)
      is deferred;
      ---Level: Public
      ---Purpose: Begins a new page of graphics in the plotter file name.

  Close (me: mutable)
--      is virtual protected;
      is virtual;
      ---C++: alias ~
      ---Level: Internal 

  Spool (me      : mutable;
      aPlotMode    : PlotMode from Aspect = Aspect_PM_FILEONLY;
      aReserved1   : CString  from Standard = NULL;
      aReserved2   : Boolean  from Standard = Standard_False)
      returns Boolean from Standard
  is virtual;
      ---Purpose:
      ---Level: Public
      
  ----------------------------------------------------------
  -- Category: Methods to create the attributes which the
  --           driver can manage itself
  ----------------------------------------------------------
  CreateDriverColorMap (me: mutable) 
  is virtual protected;
      ---Category: Methods to define standard ColorIndexs 
      ---Level: Private

  CreateDriverTypeMap (me: mutable)
  is virtual protected;
      ---Category: Methods to define standard TypeIndexs
      ---Level: Private

  CreateDriverWidthMap (me: mutable)
  is virtual protected;
      ---Category: Methods to define standard WidthIndexs
      ---Level: Private

  CreateDriverMarkMap (me: mutable)
  is virtual protected;
      ---Category: Methods to define standard MarkIndexs
      ---Level: Private

  ---------------------------------------------
  -- Category: Methods to define the attributes
  ---------------------------------------------
  InitializeColorMap (me: mutable; aColorMap: ColorMap from Aspect) 
  is virtual protected;
      ---Category: Methods to define the ColorIndexs
      ---Level: Private

  InitializeTypeMap (me: mutable; aTypeMap: TypeMap from Aspect)
  is virtual protected;
      ---Category: Methods to define the TypeIndexs
      ---Level: Private

  InitializeWidthMap (me: mutable; aWidthMap: WidthMap from Aspect)
  is virtual protected;
      ---Category: Methods to define the WidthIndexs
      ---Level: Private

  InitializeFontMap (me: mutable; aFontMap: FontMap from Aspect)
  is virtual protected;
      ---Category: Methods to define the FontIndexs
      ---Level: Private

  InitializeMarkMap (me: mutable; aFontMap: MarkMap from Aspect)
  is virtual protected;
      ---Category: Methods to define the MarkIndexs
      ---Level: Private

  ------------------------------------
  -- Methods to set graphic attributes
  ------------------------------------
  SetLineAttrib (me: mutable;
      ColorIndex: Integer from Standard;
      TypeIndex: Integer from Standard;
      WidthIndex: Integer from Standard)
  is virtual;
      ---Category: Methods to define the Current Line Attibutes
      ---Level: Public

  SetTextAttrib (me: mutable;
      ColorIndex: Integer from Standard;
      FontIndex: Integer from Standard)
  is virtual;
      ---Category: Methods to define the Current Text Attributes
      ---Level: Public

  SetTextAttrib (me: mutable;
      ColorIndex: Integer from Standard;
      FontIndex: Integer from Standard;
      aSlant: PlaneAngle from Quantity;
      aHScale: Factor from Quantity;
      aWScale: Factor from Quantity;
      isUnderlined: Boolean from Standard = Standard_False)
  is virtual;
      ---Category: Methods to define the Current Extended Text Attributes
      ---Level: Public

  SetPolyAttrib (me: mutable;
      ColorIndex: Integer from Standard;
      TileIndex: Integer from Standard;
      DrawEdge: Boolean from Standard = Standard_False)
  is virtual;
      ---Category: Methods to set the poly attributes
      ---Level: Public

  SetMarkerAttrib (me: mutable;
      ColorIndex: Integer from Standard;
      WidthIndex: Integer from Standard;
      FillMarker: Boolean from Standard = Standard_False)
  is virtual;
      ---Category: Methods to define the Current Marker Attributes
      ---Level: Public

  SetPixelSize (me: mutable ; aSize: Real from Standard)
  is static;
      ---Purpose:
      ---Level: Public

  SetPlotter (me: mutable; aPlotter: Plotter from PlotMgt)
  is static protected;
      ---Purpose: Set the plotter to be used by Spool() method.
      -- Fail if Plotter is already defined
      ---Level: Public

  --------------------------------
  -- Actual set graphic attributes
  --------------------------------
  PlotLineAttrib (me: mutable;
    ColorIndex: Integer from Standard;
    TypeIndex: Integer from Standard;
    WidthIndex: Integer from Standard)
  is virtual protected;
      ---Purpose: retrieve current line attributes
      ---Level: Private

  PlotPolyAttrib (me: mutable;
    ColorIndex: Integer from Standard;
    TileIndex: Integer from Standard;
    DrawEdge: Boolean from Standard)
  is virtual protected;
      ---Purpose: retrieve current poly attributes
      ---Level: Private

  -------------------------------------------------
  -- Incremental methods to draw graphic primitives
  -------------------------------------------------
  BeginPolyline (me : mutable; aNumber : Integer)
  is virtual;
      ---Purpose: Begin an incremental polyline primitive of <aNumber> of points .
      --  Warning: Points must be added by the the DrawPoint() method.
      ---Level: Public

  BeginPolygon (me : mutable; aNumber : Integer)
  is virtual;
      ---Purpose: Begin an incremental polygon primitive of <aNumber> of points .
      --  Warning: Points must be added by the the DrawPoint() method.
      ---Level: Public

  BeginSegments (me : mutable)
  is virtual;
      ---Purpose: Begin a set of segments.
      --  Warning: Segments must be added by the DrawSegment() method.
      ---Level: Public

  BeginArcs (me : mutable)
  is virtual;
      ---Purpose: Begin a set of circles or ellipses.
      --  Warning: Arcs must be added by the DrawArc() methods.
      ---Level: Public

  BeginPolyArcs (me : mutable)
  is virtual;
      ---Purpose: Begin a set of polygon circles or ellipses.
      --  Warning: Arcs must be added by the DrawPolyArc() methods.
      ---Level: Public

  BeginMarkers (me : mutable)
  is virtual;
      ---Purpose: Begin a set of markers.
      --  Warning: Markers must be added by the DrawMarker() method.
      ---Level: Public

  BeginPoints (me : mutable)
  is virtual;
      ---Purpose: Begin a set of points.
      --  Warning: Points must be added by the DrawPoint() method.
      ---Level: Public

  ClosePrimitive (me : mutable)
  is virtual;
      ---Purpose: Close the last Begining primitive
      ---Level: Public

  -----------------------------------------
  -- Category: Methods to manage the images
  -----------------------------------------
  IsKnownImage(me: mutable; anImage: Transient from Standard)
  returns Boolean from Standard is virtual;
      ---Purpose:
      ---Level: Public

  SizeOfImageFile (me; anImageFile: CString from Standard;
                       aWidth,aHeight: out Integer from Standard)
  returns Boolean from Standard is virtual;
      ---Purpose: Returns Standard_True and the Image Size in PIXEL
      --          if the image file exist and can be computed by the driver,
      ---Category: Methods to manage the images
      ---Level: Public

  ClearImage (me: mutable; anImageId: Transient from Standard)
  is virtual;
      ---Purpose:
      ---Level: Public

  ClearImageFile (me: mutable; anImageFile: CString from Standard)
  is virtual;
      ---Purpose: Clears the image associated with the image file .
      ---Category: Methods to manage the images
      ---Level: Public

  DrawImage (me: mutable; anImageId: Transient from Standard;
             aX, aY: ShortReal from Standard)
  is virtual;
      ---Purpose: Draws the image  in <me>.
      --          <aX>, <aY> is the center of the image.
      --          Image center must be defined in DPU space.
      ---Category: Methods to manage the images
      ---Level: Public

  DrawImageFile (me: mutable; anImageFile: CString from Standard;
                 aX, aY: ShortReal from Standard;
                 aScale: Factor from Quantity = 1.0)
  is virtual;
      ---Purpose: Draws the image file in <me>.
      --          <aX>, <aY> is the center of the image.
      --          Image center must be defined in DPU space.
      ---Category: Methods to manage the images
      ---Level: Public
  
  FillAndDrawImage (me: mutable; anImageId: Transient from Standard;
      aX, aY: ShortReal from Standard;
      aWidth, aHeight: Integer from Standard;
      anArrayOfPixels: Address from Standard)
  is virtual;
      ---Purpose: Draw a complete image .
      --          Image size must be defined in DPU space>
      ---Category: Methods to manage the images
      ---Level: Public
 

  FillAndDrawImage (me: mutable; anImageId: Transient from Standard;
      aX, aY: ShortReal from Standard;
      anIndexOfLine, aWidth, aHeight: Integer from Standard;
      anArrayOfPixels: Address from Standard)
  is virtual;
      ---Purpose: Fills a line of the Image .
      ---Category: Methods to manage the images
      ---Level: Public

  -------------------------------------
  -- Methods to draw graphic primitives
  -------------------------------------
  DrawPoint (me : mutable; X, Y: ShortReal from Standard)
  is static;
      ---Purpose: Draws a 1 PIXEL point depending of the SetMarkerAttrib()
      --color attribute or add a point depending of the incremental BeginXxxxxx()
      --primitive used.
      ---Category: Methods to draw primitives
      ---Level: Public


  DrawSegment (me : mutable;
      X1, Y1: ShortReal from Standard;
      X2, Y2: ShortReal from Standard)
  is static;
      ---Purpose: Draw a segment depending of the SetLineAttrib() attributes.
      ---Category: Methods to draw primitives
      ---Level: Public


  DrawRectangle (me : mutable; aX,aY : ShortReal from Standard;
      aDX,aDY : ShortReal from Standard)
  is static;
      ---Purpose: Draw a rectangle. aX,aY is start point
      --      aDX , aDY are horizontal and vertical dimensions
      ---Level: Public


  DrawPolyline (me : mutable;
      aListX, aListY: Array1OfShortReal from TShort)
  is static;
      ---Purpose: Draw a polyline depending of the SetLineAttrib() attributes.
      ---Category: Methods to draw primitives
      ---Level: Public


  DrawPolygon (me : mutable;
      aListX, aListY: Array1OfShortReal from TShort)
  is static;
      ---Purpose: Draw a polygon depending of the SetPolyAttrib() attributes. 
      ---Category: Methods to draw primitives
      ---Level: Public


  DrawArc (me : mutable; X,Y : ShortReal from Standard;
      anXradius,anYradius : ShortReal from Standard;
      aStartAngle: ShortReal from Standard = 0.0;
      anOpenAngle: ShortReal from Standard = 6.283185) 
  returns Boolean from Standard
  is static;
      ---Purpose: Draws an Ellipsoid arc of center <X,Y> and Radius
      --<anXradius,anYradius> of relative angle <anOpenAngle> from 
      --the base angle <aStartAngle> and depending of the SetLineAttrib() attributes.
      --  Warning: Returns FALSE if the hardware can't drawing this
      --primitive properly,application must to simulate it.        
      ---Category: Methods to draw primitives
      ---Level: 


  DrawPolyArc (me : mutable; X,Y : ShortReal from Standard;
      anXradius,anYradius : ShortReal from Standard;
      aStartAngle: ShortReal from Standard = 0.0;
      anOpenAngle: ShortReal from Standard = 6.283185)
  returns Boolean from Standard
  is static;
      ---Purpose: Draws an filled Ellipsoid arc of center <X,Y> and Radius
      --<anXradius,anYradius> of relative angle <anOpenAngle> from 
      --the base angle <aStartAngle> and depending of the SetPolyAttrib() attributes.
      --  Warning: Returns FALSE if the hardware can't drawing this
      --primitive properly,application must to simulate it.           
      ---Category: Methods to draw primitives
      ---Level: Public


  DrawMarker (me : mutable;
      aMarker: Integer from Standard;
      Xpos:  ShortReal from Standard;
      Ypos:  ShortReal from Standard;
      Width: ShortReal from Standard;
      Height: ShortReal from Standard;
      Angle: ShortReal from Standard = 0.0)
  is static;
      ---Purpose: Draws the marker <aMarker>
      --depending of the SetMarkerAttrib() attributes.
      --  Warning: Coordinates and sizes must be defined in DWU space.
      --      Angle must be defined in RADIAN.
      --      A one pixel marker is drawn when aMarker index is undefined.
      ---Category: Methods to draw primitives
      ---Level: Public


  DrawText (me : mutable;
      aText: ExtendedString from TCollection;
      Xpos:  ShortReal from Standard;
      Ypos:  ShortReal from Standard;
      anAngle: ShortReal from Standard = 0.0;
      aType: TypeOfText from Aspect = Aspect_TOT_SOLID)
  is static;
      ---Purpose: Draws a text depending of the SetTextAttrib() attributes.
      --  Warning: Coordinates must be defined in DWU space.
      ---Category: Methods to draw primitives
      ---Level: Public


  DrawText (me : mutable;
      aText: CString from Standard;
      Xpos:  ShortReal from Standard;
      Ypos:  ShortReal from Standard;
      anAngle: ShortReal from Standard = 0.0;
      aType: TypeOfText from Aspect = Aspect_TOT_SOLID)
  is static;
      ---Purpose: Draws a text depending of the SetTextAttrib() attributes.
      --  Warning: Coordinates must be defined in DWU space.
      ---Category: Methods to draw primitives
      ---Level: Public


  DrawPolyText (me : mutable;
      aText: ExtendedString from TCollection;
      Xpos:  ShortReal from Standard;
      Ypos:  ShortReal from Standard;
      aMargin: Ratio from Quantity = 0.1;
      anAngle: ShortReal from Standard = 0.0;
      aType: TypeOfText from Aspect = Aspect_TOT_SOLID)
  is static;
      ---Purpose: Draws an framed text depending of the
      -- SetTextAttrib() and SetPolyAttrib() attributes.
      --  Warning: Coordinates must be defined in DWU space.
      --          <aMarge> defines the ratio of the space between the
      --          polygon borders and the bounding box of the text and
      --          depending of the height of the text.
      ---Category: Methods to draw primitives
      ---Level: Public


  DrawPolyText (me : mutable;
      aText: CString from Standard;
      Xpos:  ShortReal from Standard;
      Ypos:  ShortReal from Standard;
      aMargin: Ratio from Quantity = 0.1;
      anAngle: ShortReal from Standard = 0.0;
      aType: TypeOfText from Aspect = Aspect_TOT_SOLID)
  is static;
      ---Purpose: Draws an framed text depending of the
      -- SetTextAttrib() and SetPolyAttrib() attributes.
      --  Warning: Coordinates must be defined in DWU space.
      --          <aMarge> defines the ratio of the space between the
      --          polygon borders and the bounding box of the text and
      --          depending of the height of the text.
      ---Category: Methods to draw primitives
      ---Level: Public


  --------------------------------------------------
  -- Private plot methods to draw graphic primitives
  --------------------------------------------------
  PlotPoint (me : mutable; X, Y: ShortReal from Standard)
  returns Boolean from Standard
  is virtual protected;
      ---Purpose:
      ---Category:
      ---Level: Private


  PlotSegment (me : mutable;
      X1, Y1: ShortReal from Standard;
      X2, Y2: ShortReal from Standard)
  returns Boolean from Standard
  is virtual protected;
      ---Purpose:
      ---Category:
      ---Level: Private


  PlotRectangle (me : mutable; aX,aY : ShortReal from Standard;
      aDX,aDY : ShortReal from Standard;
      aAngle: ShortReal from Standard = 0.0)
  returns Boolean        
  is virtual protected;
      ---Purpose:
      ---Category:
      ---Level: Private


  PlotPolyline (me : mutable;
      xArray : Address from Standard;
      yArray : Address from Standard;
      nPts   : Address from Standard;
      nParts : Integer from Standard)
  returns Boolean from Standard
  is virtual protected;
      ---Purpose:
      ---Category:
      ---Level: Private


  PlotPolygon (me : mutable;
      xArray : Address from Standard;
      yArray : Address from Standard;
      nPts   : Address from Standard;
      nParts : Integer from Standard)
  returns Boolean from Standard
  is virtual protected;
      ---Purpose:
      ---Category:
      ---Level: Private


  PlotArc (me : mutable; X,Y : ShortReal from Standard;
      anXradius,anYradius : ShortReal from Standard;
      sAngle: ShortReal from Standard;
      oAngle: ShortReal from Standard)
  returns Boolean from Standard
  is virtual protected;
      ---Purpose:
      ---Category:
      ---Level: Private


  PlotPolyArc (me : mutable; X,Y : ShortReal from Standard;
      anXradius,anYradius : ShortReal from Standard;
      sAngle: ShortReal from Standard;
      oAngle: ShortReal from Standard)
  returns Boolean from Standard
  is virtual protected;
      ---Purpose:
      ---Category:
      ---Level: Private


  PlotMarker (me : mutable;
      aMarker: Integer from Standard;
      Xpos:  ShortReal from Standard;
      Ypos:  ShortReal from Standard;
      Width: ShortReal from Standard;
      Height: ShortReal from Standard;
      Angle: ShortReal from Standard)
  returns Boolean from Standard
  is virtual protected;
      ---Purpose:
      ---Category:
      ---Level: Private


  PlotText (me : mutable;
      aText: ExtendedString from TCollection;
      Xpos:  ShortReal from Standard;
      Ypos:  ShortReal from Standard;
      anAngle: ShortReal from Standard;
      aType: TypeOfText from Aspect)
  returns Boolean from Standard
  is virtual protected;
      ---Purpose:
      ---Category:
      ---Level: Private
      

  PlotText (me : mutable;
      aText: CString from Standard;
      Xpos:  ShortReal from Standard;
      Ypos:  ShortReal from Standard;
      anAngle: ShortReal from Standard;
      aType: TypeOfText from Aspect)
  returns Boolean from Standard
  is virtual protected;
      ---Purpose:
      ---Category:
      ---Level: Private


  PlotPolyText (me : mutable;
      aText: ExtendedString from TCollection;
      Xpos:  ShortReal from Standard;
      Ypos:  ShortReal from Standard;
      aMargin: Ratio from Quantity;
      anAngle: ShortReal from Standard;
      aType: TypeOfText from Aspect)
  returns Boolean from Standard
  is virtual protected;
      ---Purpose:
      ---Category:
      ---Level: Private


  PlotPolyText (me : mutable;
      aText: CString from Standard;
      Xpos:  ShortReal from Standard;
      Ypos:  ShortReal from Standard;
      aMargin: Ratio from Quantity;
      anAngle: ShortReal from Standard;
      aType: TypeOfText from Aspect)
  returns Boolean from Standard
  is virtual protected;
      ---Purpose:
      ---Category:
      ---Level: Private


  PlotImage (me: mutable; 
      aX, aY, aWidth:  ShortReal from Standard;
      aHeight, aScale: ShortReal from Standard;
      anImageFile:     CString   from Standard;
      anArrayOfPixels: Address   from Standard;
      aLineIndex:      Integer   from Standard = -1)
  returns Boolean from Standard
  is virtual protected;
      ---Purpose:
      ---Category:
      ---Level: Private


  ----------------------------------------------------
  --- Inquire methods
  ----------------------------------------------------
  Plotter (me)
    returns Plotter from PlotMgt;
      ---Purpose:
      ---Category: Inquire methods
      ---Level: Public

  Cout (me)
    returns FStream from Aspect
    is static protected;
      ---Purpose:
      ---Category: Inquire methods
      ---Level: Public

  PlotFileName (me)
    returns AsciiString from TCollection;
      ---Purpose:
      ---Category: Inquire methods
      ---Level: Public

  DrawingName (me)
    returns AsciiString from TCollection;
      ---Purpose:
      ---Category: Inquire methods
      ---Level: Public

  SpoolDirectory (me)
    returns AsciiString from TCollection;
      ---Purpose:
      ---Category: Inquire methods
      ---Level: Public

  WorkSpace (me ; Width,Height : out Length from Quantity)
  is redefined;
      ---Purpose: Returns the Available WorkSpace in DWU coordinates
      ---Category: Inquire methods
      ---Level: Public

  Convert (me; PV : Integer from Standard)
    returns Length from Quantity is redefined virtual;
      ---Purpose: Returns the DWU value depending of the PIXEL value.
      ---Category: Inquire methods
      ---Level: Public

  Convert (me; DV : Length from Quantity)
    returns Integer from Standard is redefined virtual;
      ---Purpose: Returns the PIXEL value depending of the DWU value.
      ---Category: Inquire methods
      ---Level: Public

  Convert (me; PX, PY : Integer from Standard;
      DX, DY : out Length from Quantity) is redefined virtual;
      ---Purpose: Returns the DWU position depending of the PIXEL position.
      ---Category: Inquire methods
      ---Level: Public

  Convert (me; DX, DY : Length from Quantity;
      PX, PY : out Integer from Standard) is redefined virtual;
      ---Purpose: Returns the PIXEL position depending of the DWU position .
      ---Category: Inquire methods
      ---Level: Public

  LineAttrib (me; ColorIndex, TypeIndex, WidthIndex : out Integer from Standard);
      ---Purpose:
      ---Category: Inquire methods
      ---Level: Public

  PolyAttrib (me; ColorIndex, TileIndex : out Integer from Standard;
                  EdgeFlag : out Boolean from Standard);
      ---Purpose:
      ---Category: Inquire methods
      ---Level: Public

  DrawCurveCapable (me)
  returns Boolean from Standard is virtual protected;
      ---Purpose: Should be called from PlotMgt_TextManager::Curveto()
      ---         method to check if the driver is capable to draw curves.
      ---Category: Inquire methods
      ---Level: Private

  MapX(me; aShortReal: ShortReal from Standard) 
  returns ShortReal from Standard is virtual private;
      ---Purpose:
      ---Category: Inquire methods
      ---Level: Private

  MapY(me; aShortReal: ShortReal from Standard) 
  returns ShortReal from Standard is virtual private;
      ---Purpose:
      ---Category: Inquire methods
      ---Level: Private

fields
  myFStream          : FStream           from Aspect;
  myPixelSize        : Real              from Standard is protected;
  myDrawingName      : AsciiString       from TCollection is protected;
  myFileName         : AsciiString       from TCollection is protected;
  myPlotter          : Plotter           from PlotMgt;
  myPlotterIsDefined : Boolean           from Standard;

  ----- Draw attibutes
  myWidth            : ShortReal         from Standard is protected;
  myHeight           : ShortReal         from Standard is protected;
  myPaperMargin      : ShortReal         from Standard is protected;
  myTypeOfColorSpace : TypeOfColorSpace  from Aspect is protected;

  ----- Actual attributes (written in the file)
  myColorIndex       : Integer           from Standard is protected;
  myTypeIndex        : Integer           from Standard is protected;
  myWidthIndex       : Integer           from Standard is protected;
  myFontIndex        : Integer           from Standard is protected;

  ----- Graphic attributes (set by SetXXX methods)
  myLineColorIndex   : Integer           from Standard is protected;
  myLineTypeIndex    : Integer           from Standard is protected;
  myLineWidthIndex   : Integer           from Standard is protected;

  myPolyColorIndex   : Integer           from Standard is protected;
  myPolyTileIndex    : Integer           from Standard is protected;
  myPolyEdgeFlag     : Boolean           from Standard is protected;

  myMarkerColorIndex : Integer           from Standard is protected;
  myMarkerWidthIndex : Integer           from Standard is protected;
  myMarkerFillFlag   : Boolean           from Standard is protected;

  myTextColorIndex   : Integer           from Standard is protected;
  myTextFontIndex    : Integer           from Standard is protected;
  myTextHScale       : Real              from Standard is protected;
  myTextWScale       : Real              from Standard is protected;
  myTextSlant        : Real              from Standard is protected;
  myTextMinHeight    : Real              from Standard is protected;
  myTextIsUnderlined : Boolean           from Standard is protected;
  myCapsHeight       : Boolean           from Standard is protected;

  ----- Interal attributes and parameters
  myPrimitiveType    : TypeOfPrimitive   from Aspect is protected;
  myPrimitiveLength  : Integer           from Standard is protected;
  myPrimitiveX       : Array1OfShortReal from TShort is protected;
  myPrimitiveY       : Array1OfShortReal from TShort is protected;

  myMFTFonts         : HListOfMFTFonts   from PlotMgt is protected;
  myMFTSizes         : HArray1OfShortReal from TShort is protected;
  myTextManager      : TextManager       from PlotMgt is protected;

  ----- Private attributes, supported by the driver
  myDriverColorMap   : ColorMap          from Aspect is protected;
  myDriverTypeMap    : TypeMap           from Aspect is protected;
  myDriverWidthMap   : WidthMap          from Aspect is protected;
  myDriverMarkMap    : MarkMap           from Aspect is protected;
  
friends
  class TextManager from PlotMgt

end PlotterDriver from PlotMgt;
