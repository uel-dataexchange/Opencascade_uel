-- File:	MakeElips.cdl
-- Created:	Wed Aug 26 14:31:40 1992
-- Author:	Remi GILET
--		<reg@topsn3>
---Copyright:	 Matra Datavision 1992

class MakeElips from gce inherits Root from gce

    	---Purpose :This class implements the following algorithms used to 
    	--          create an ellipse from gp.
    	--          
    	--          * Create an ellipse from its center, and two points:
    	--            one on the ciconference giving the major radius, the 
    	--            other giving the value of the small radius.

uses Pnt   from gp,
     Ax2   from gp,
     Elips from gp

raises NotDone from StdFail

is

Create (A2 :                       Ax2  from gp;
        MajorRadius, MinorRadius : Real from Standard) 
    returns MakeElips;
    	--- Purpose :The major radius of the ellipse is on the "XAxis" and the
    	--           minor radius is on the "YAxis" of the ellipse. The "XAxis"
    	--           is defined with the "XDirection" of A2 and the "YAxis" is
    	--           defined with the "YDirection" of A2.
    	-- Warnings :
    	--           It is not forbidden to create an ellipse with 
    	--           MajorRadius = MinorRadius.

Create(S1,S2  : Pnt from gp;
       Center : Pnt from gp) returns MakeElips;
	---Purpose: Make an ellipse with its center and two points.
	-- Warning
    	-- The MakeElips class does not prevent the
    	-- construction of an ellipse where the MajorRadius is
    	-- equal to the MinorRadius.
    	-- If an error occurs (that is, when IsDone returns
    	-- false), the Status function returns:
    	-- -   gce_InvertRadius if MajorRadius is less than MinorRadius;
    	-- -   gce_NegativeRadius if MinorRadius is less than 0.0;
    	-- -   gce_NullAxis if the points S1 and Center are coincident; or
    	-- -   gce_InvertAxis if:
    	--   -   the major radius computed with Center and S1
    	--    is less than the minor radius computed with Center, S1 and S2, or
    	--   -   Center, S1 and S2 are collinear.         
		
Value(me) returns Elips from gp
    raises NotDone
    is static;
      	---C++: return const&
    	---Purpose: Returns the constructed ellipse.
    	-- Exceptions StdFail_NotDone if no ellipse is constructed.   
    
Operator(me) returns Elips from gp
    is static;
    	---C++: return const&
    	---C++: alias "Standard_EXPORT operator gp_Elips() const;"

fields

    TheElips : Elips from gp;
    --The solution from gp.
    
end MakeElips;




