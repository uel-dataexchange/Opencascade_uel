-- File:	BRepAlgoAPI_Fuse.cdl
-- Created:	Thu Oct 14 18:24:07 1993
-- Author:	Remi LEQUETTE
--		<rle@phylox>
---Copyright:	 Matra Datavision 1993



class Fuse from BRepAlgoAPI inherits BooleanOperation from BRepAlgoAPI

	---Purpose:  The class Fuse provides a
    	-- Boolean fusion operation on a pair of arguments (Boolean Union).
    	-- The class Fuse provides a framework for:
    	--   -       Defining the construction of a fused shape;
    	--   -       Implementing the building algorithm
    	--   -       Consulting the result.

uses
    Shape from TopoDS, 
    DSFiller from BOPTools

is
    Create (S1,S2 : Shape from TopoDS)  
    	returns Fuse from BRepAlgoAPI;  
	---Purpose: Constructs a fuse of shapes aS1 and aS2.
	 
    Create (S1,S2 : Shape from TopoDS; 
    	    aDSF:DSFiller from BOPTools)  
    	returns Fuse from BRepAlgoAPI; 
    
    	---Purpose: Constructs a new shape that is a fuse of shapes aS1 and aS2 using aDSFiller. 
    
end Fuse;
