-- File:	IGESGraph_ToolPick.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolPick  from IGESGraph

    ---Purpose : Tool to work on a Pick. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses Pick from IGESGraph,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolPick;
    ---Purpose : Returns a ToolPick, ready to work


    ReadOwnParams (me; ent : mutable Pick;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : Pick;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : Pick;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a Pick <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable Pick) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a Pick
    --           (NbPropertyValues forced to 1)

    DirChecker (me; ent : Pick) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : Pick;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : Pick; entto : mutable Pick;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : Pick;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolPick;
