-- File:	StepToGeom_MakeCurve2d.cdl
-- Created:	Wed Aug  4 10:42:37 1993
-- Author:	Martine LANGLOIS
---Copyright:	 Matra Datavision 1993

class MakeCurve2d from StepToGeom

    ---Purpose: This class implements the mapping between 
    --          class Curve from StepGeom which
    --          describes a Curve from prostep and Curve from Geom2d. 
    --          As Curve is an abstract class
    --          this class an access to the sub-class required.

uses Curve from Geom2d,
     Curve from StepGeom

is 

    Convert ( myclass; SC : Curve from StepGeom;
                       CC : out Curve from Geom2d )
    returns Boolean from Standard;

end MakeCurve2d;
