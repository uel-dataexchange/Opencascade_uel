--
-- Package: OpenGl
-- Author:  CAL
-- Created: Mercredi 4 Janvier 1995
-- Updated: 20/08/97 ; PCT : ajout texture mapping
--      27/01/98 ; FMN : Delete GEOMLITE
--              
-- Copyright:   MatraDatavision 1995
--
-- Purpose: Specifications definitives
--

package OpenGl

    ---Version:

    ---Purpose: This package contains the common OpenGl graphic interface.

    ---Keywords: OpenGl, CInterface

    ---Warning: No class in this package. It is used only to archive
    --      all the objects files in a library.
    ---References:

uses

    OSD,
    TColStd,
    TCollection,
    Aspect,
    Quantity,
    Graphic3d,
    Image, 
    AlienImage

is

    exception Error inherits NumericError from Standard;

    class GraphicDriver;
    ---Purpose: Defines a graphic driver for the opengl interface

end OpenGl;
