-- File:	IGESDraw_ToolCircArraySubfigure.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolCircArraySubfigure  from IGESDraw

    ---Purpose : Tool to work on a CircArraySubfigure. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses CircArraySubfigure from IGESDraw,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolCircArraySubfigure;
    ---Purpose : Returns a ToolCircArraySubfigure, ready to work


    ReadOwnParams (me; ent : mutable CircArraySubfigure;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : CircArraySubfigure;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : CircArraySubfigure;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a CircArraySubfigure <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : CircArraySubfigure) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : CircArraySubfigure;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : CircArraySubfigure; entto : mutable CircArraySubfigure;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : CircArraySubfigure;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolCircArraySubfigure;
