-- File:	ShapeUpgrade_ShapeDivideClosed.cdl
-- Created:	Thu Jul 22 17:58:21 1999
-- Author:	data exchange team
--		<det@friendox>
---Copyright:	 Matra Datavision 1999


class ShapeDivideClosed from ShapeUpgrade inherits ShapeDivide from ShapeUpgrade

	---Purpose: Divides all closed faces in the shape. Class 
    	--          ShapeUpgrade_ClosedFaceDivide is used as divide tool.

uses

    Shape from TopoDS

is
    Create (S: Shape from TopoDS) returns ShapeDivideClosed from ShapeUpgrade;
    	---Purpose: Initialises tool with shape and default parameter.
    
    SetNbSplitPoints (me: in out; num: Integer);
    	---Purpose: Sets the number of cuts applied to divide closed faces.
	--          The number of resulting faces will be num+1.
    

end ShapeDivideClosed;
