-- File:	Transfer_BinderOfTransientInteger.cdl
-- Created:	Mon Feb 27 15:06:40 1995
-- Author:	Christian CAILLET
--		<cky@anion>
---Copyright:	 Matra Datavision 1995


class BinderOfTransientInteger  from Transfer  inherits SimpleBinderOfTransient

    ---Purpose : This type of Binder allows to attach as result, besides a
    --           Transient Object, an Integer Value, which can be an Index
    --           in the Object if it defines a List, for instance
    --           
    --           This Binder is otherwise a kind of SimpleBinderOfTransient,
    --           i.e. its basic result (for iterators, etc) is the Transient

uses Integer

is

    Create returns mutable BinderOfTransientInteger;
    ---Purpose : Creates an empty BinderOfTransientInteger; Default value for
    --           the integer part is zero

    SetInteger (me : mutable; value : Integer);
    ---Purpose : Sets a value for the integer part

    Integer (me) returns Integer;
    ---Purpose : Returns the value set for the integer part

fields

    theintval : Integer;

end BinderOfTransientInteger;
