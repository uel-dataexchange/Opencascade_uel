-- File:	IGESSelect_SelectBypassSubfigure.cdl
-- Created:	Tue Jan 13 08:44:11 1998
-- Author:	Christian CAILLET
--		<xstep@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1998


class SelectBypassSubfigure  from IGESSelect  inherits SelectExplore

    ---Purpose : Selects a list built as follows :
    --           Subfigures correspond to
    --           * Definition (basic : type 308, or Network : type 320)
    --           * Instance (Singular : type 408, or Network : 420, or
    --             patterns : 412,414)
    --           
    --           Entities which are not Subfigure are taken as such
    --           For Subfigures Instances, their definition is taken, then
    --           explored itself
    --           For Subfigures Definitions, the list of "Associated Entities"
    --           is explored
    --           Hence, level 0 (D) recursively explores a Subfigure if some of
    --           its Elements are Subfigures. level 1 explores just at first
    --           level (i.e. for an instance, returns its definition)

uses AsciiString from TCollection, Transient, EntityIterator, Graph

raises InterfaceError

is

    Create (level : Integer = 0) returns mutable SelectBypassSubfigure;
    ---Purpose : Creates a SelectBypassSubfigure, by default all level
    --           (level = 1 explores at first level)

    Explore (me; level : Integer; ent : Transient; G : Graph;
    	     explored : in out EntityIterator)
    	returns Boolean;
    ---Purpose : Explores an entity : for a Subfigure, gives its elements
    --           Else, takes the entity itself


    ExploreLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium : "Content of Subfigure"

end SelectBypassSubfigure;
