-- File:        Address.cdl
-- Created:     Mon Dec  4 12:02:22 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWAddress from RWStepBasic

	---Purpose : Read & Write Module for Address

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Address from StepBasic

is

	Create returns RWAddress;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Address from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : Address from StepBasic);

end RWAddress;
