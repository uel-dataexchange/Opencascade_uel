-- File:        Axis2Placement2d.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWAxis2Placement2d from RWStepGeom

	---Purpose : Read & Write Module for Axis2Placement2d

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Axis2Placement2d from StepGeom,
     EntityIterator from Interface

is

	Create returns RWAxis2Placement2d;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Axis2Placement2d from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : Axis2Placement2d from StepGeom);

	Share(me; ent : Axis2Placement2d from StepGeom; iter : in out EntityIterator);

end RWAxis2Placement2d;
