-- File:	RWStepBasic_RWDocumentFile.cdl
-- Created:	Thu May 11 16:38:00 2000 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWDocumentFile from RWStepBasic

    ---Purpose: Read & Write tool for DocumentFile

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    DocumentFile from StepBasic

is
    Create returns RWDocumentFile from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : DocumentFile from StepBasic);
	---Purpose: Reads DocumentFile

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: DocumentFile from StepBasic);
	---Purpose: Writes DocumentFile

    Share (me; ent : DocumentFile from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWDocumentFile;
