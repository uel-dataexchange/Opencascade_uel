-- File:        RepresentationContext.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWRepresentationContext from RWStepRepr

	---Purpose : Read & Write Module for RepresentationContext

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     RepresentationContext from StepRepr

is

	Create returns RWRepresentationContext;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable RepresentationContext from StepRepr);

	WriteStep (me; SW : in out StepWriter; ent : RepresentationContext from StepRepr);

end RWRepresentationContext;
