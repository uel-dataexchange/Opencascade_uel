-- File:	LocOpe_ProjectedWires.cdl
-- Created:	Mon Jan  8 16:03:41 1996
-- Author:	Jacques GOUSSARD
--		<jag@bravox>
---Copyright:	 Matra Datavision 1996


deferred class ProjectedWires from LocOpe inherits TShared from MMgt

	---Purpose: 

uses Face   from TopoDS,
     Wire   from TopoDS,
     Edge   from TopoDS,
     Vertex from TopoDS

is

    InitEdgeIterator(me: mutable)
    
    	is deferred;


    MoreEdge(me: mutable)
    	returns Boolean from Standard
	is deferred;


    Edge(me: mutable)
    	returns Edge from TopoDS
	is deferred;


    OnFace(me: mutable)
	---Purpose: Returns the face of the shape on which the current
	--          edge is projected.
    	returns Face from TopoDS
	is deferred;

    
    OnEdge(me: mutable; E: out Edge from TopoDS)
	---Purpose: If the   current  edge is  projected  on  an edge,
	--          returns <Standard_True> and sets the value of <E>.
	--          Otherwise, returns <Standard_False>.
    	returns Boolean from Standard
	is deferred;


    NextEdge(me: mutable)
    
    	is deferred;


    OnVertex(me: mutable; Vwire :     Vertex from TopoDS;
    	                  Vshape: out Vertex from TopoDS)
			  
	returns Boolean from Standard
	is deferred;


    OnEdge(me: mutable; V: Vertex from TopoDS;
                        E: out Edge from TopoDS;
			P: out Real from Standard)
	---Purpose: If the vertex <V> lies on  an edge of the original
	--          shape,  returns     <Standard_True> and   sets the
	--          concerned edge in  <E>,  and the parameter on  the
	--          edge in <P>.
	--          Else returns <Standard_False>.
	returns Boolean from Standard
	is deferred;


end ProjectedWires;
