-- File:	StepAP214_AppliedPersonAndOrganizationAssignment.cdl
-- Created:	Tue Mar  9 15:29:30 1999
-- Author:	data exchange team
--		<det@androx.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class AppliedPersonAndOrganizationAssignment from StepAP214 

inherits PersonAndOrganizationAssignment from StepBasic
       

uses
    
    	HArray1OfPersonAndOrganizationItem from StepAP214,
    	PersonAndOrganizationItem from StepAP214,
    	PersonAndOrganization from StepBasic,
    	PersonAndOrganizationRole from StepBasic

is
    	Create returns mutable AppliedPersonAndOrganizationAssignment;
	---Purpose: Returns a AutoDesignDateAndPersonAssignment
	
	Init (me : mutable;
	      aAssignedPersonAndOrganization : mutable PersonAndOrganization from StepBasic;
	      aRole : mutable PersonAndOrganizationRole from StepBasic) is redefined;
	
	Init (me : mutable;
	      aAssignedPersonAndOrganization : mutable PersonAndOrganization from StepBasic;
	      aRole : mutable PersonAndOrganizationRole from StepBasic;
	      aItems : mutable HArray1OfPersonAndOrganizationItem from StepAP214) is virtual;
	
    	-- Specific Methods for Field Data Access --
	
	SetItems(me : mutable; aItems : mutable HArray1OfPersonAndOrganizationItem);
	Items (me) returns mutable HArray1OfPersonAndOrganizationItem;
	ItemsValue (me; num : Integer) returns PersonAndOrganizationItem;
	NbItems (me) returns Integer;
	
	
fields
    items : HArray1OfPersonAndOrganizationItem from StepAP214; -- a SelectType
    
end AppliedPersonAndOrganizationAssignment;
