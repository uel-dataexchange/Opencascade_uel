-- File:	RWStepShape_RWShapeDefinitionRepresentation.cdl
-- Created:	Fri Nov 26 16:26:39 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWShapeDefinitionRepresentation from RWStepShape

    ---Purpose: Read & Write tool for ShapeDefinitionRepresentation

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ShapeDefinitionRepresentation from StepShape

is
    Create returns RWShapeDefinitionRepresentation from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ShapeDefinitionRepresentation from StepShape);
	---Purpose: Reads ShapeDefinitionRepresentation

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ShapeDefinitionRepresentation from StepShape);
	---Purpose: Writes ShapeDefinitionRepresentation

    Share (me; ent : ShapeDefinitionRepresentation from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)


end RWShapeDefinitionRepresentation;
