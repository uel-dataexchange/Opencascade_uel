-- File:	RWStepFEA_RWCurveElementEndRelease.cdl
-- Created:	Thu Dec 12 17:51:04 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWCurveElementEndRelease from RWStepFEA

    ---Purpose: Read & Write tool for CurveElementEndRelease

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    CurveElementEndRelease from StepFEA

is
    Create returns RWCurveElementEndRelease from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : CurveElementEndRelease from StepFEA);
	---Purpose: Reads CurveElementEndRelease

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: CurveElementEndRelease from StepFEA);
	---Purpose: Writes CurveElementEndRelease

    Share (me; ent : CurveElementEndRelease from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWCurveElementEndRelease;
