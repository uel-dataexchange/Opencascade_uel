-- File:	IGESSelect_RebuildGroups.cdl
-- Created:	Wed Jun  1 18:08:58 1994
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1994


class RebuildGroups  from IGESSelect  inherits ModelModifier from IGESSelect

    ---Purpose : Rebuilds Groups which were bypassed to produce new models.
    --           If a set of entities, all put into a same IGESModel, were
    --           part of a same Group in the starting Model, this Modifier
    --           rebuilds the original group, but only with the transferred
    --           entities. The distinctions (Ordered or not, "WhithoutBackP"
    --           or not) are renewed, also the name of the group.
    --           
    --           If the Input Selection is present, tries to rebuild groups
    --           only for the selected entities. Else, tries to rebuild
    --           groups for all the transferred entities.

uses AsciiString from TCollection,
     IGESModel, CopyTool, ContextModif

is

    Create returns mutable RebuildGroups;
    ---Purpose : Creates an RebuildGroups, which uses the system Date

    Performing (me; ctx : in out ContextModif;
    	        target  : mutable IGESModel;
                TC      : in out CopyTool);
    ---Purpose : Specific action : Rebuilds the original groups

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text which is
    --           "Rebuild Groups"

end RebuildGroups;
