-- File:        Sphere.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSphere from RWStepShape

	---Purpose : Read & Write Module for Sphere

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Sphere from StepShape,
     EntityIterator from Interface

is

	Create returns RWSphere;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Sphere from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : Sphere from StepShape);

	Share(me; ent : Sphere from StepShape; iter : in out EntityIterator);

end RWSphere;
