-- File:	Prs3d_LengthPresentation.cdl
-- Created:	Thu Jun  3 09:41:39 1993
-- Author:	Jean-Louis FRENKEL
--		<jlf@stylox>
---Copyright:	 Matra Datavision 1993



class LengthPresentation from Prs3d inherits Root from Prs3d
    	---Purpose: A framework to define the display of lengths.
uses
    Presentation from Prs3d,
    Pnt from gp,
    Drawer from Prs3d,
    ExtendedString from TCollection
    	
is  
    Draw( myclass; aPresentation: Presentation from Prs3d;
    	    	   aDrawer: Drawer from Prs3d;
		   aText: ExtendedString from TCollection;
                   AttachmentPoint1: Pnt from gp;
		   AttachmentPoint2: Pnt from gp;
		   OffsetPoint: Pnt from gp);
    	---Purpose: Defines the display of the length between the points
    	-- AttachmentPoint1 and AttachmentPoint2.
    	-- The text aText is displayed at the point OffsetPoint,
    	-- and the drawer aDrawer specifies the display
    	-- attributes which lengths will have.
    	-- The presentation object aPresentation stores the
    	-- information defined in this framework.
end LengthPresentation from Prs3d;
