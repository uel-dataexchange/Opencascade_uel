-- File:	RWStepBasic_RWMechanicalContext.cdl
-- Created:	Wed Jul 24 14:36:23 1996
-- Author:	Frederic MAUPAS
--		<fma@pronox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996

class RWMechanicalContext from RWStepBasic

	---Purpose : Read & Write Module for MechanicalContext

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     MechanicalContext from StepBasic,
     EntityIterator from Interface

is

	Create returns RWMechanicalContext;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable MechanicalContext from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : MechanicalContext from StepBasic);

	Share(me; ent : MechanicalContext from StepBasic; iter : in out EntityIterator);

end RWMechanicalContext;
