-- File:	StepRepr_MakeFromUsageOption.cdl
-- Created:	Mon Jul  3 20:13:36 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class MakeFromUsageOption from StepRepr
inherits ProductDefinitionUsage from StepRepr

    ---Purpose: Representation of STEP entity MakeFromUsageOption

uses
    HAsciiString from TCollection,
    ProductDefinition from StepBasic,
    MeasureWithUnit from StepBasic

is
    Create returns MakeFromUsageOption from StepRepr;
	---Purpose: Empty constructor

    Init (me: mutable; aProductDefinitionRelationship_Id: HAsciiString from TCollection;
                       aProductDefinitionRelationship_Name: HAsciiString from TCollection;
                       hasProductDefinitionRelationship_Description: Boolean;
                       aProductDefinitionRelationship_Description: HAsciiString from TCollection;
                       aProductDefinitionRelationship_RelatingProductDefinition: ProductDefinition from StepBasic;
                       aProductDefinitionRelationship_RelatedProductDefinition: ProductDefinition from StepBasic;
                       aRanking: Integer;
                       aRankingRationale: HAsciiString from TCollection;
                       aQuantity: MeasureWithUnit from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Ranking (me) returns Integer;
	---Purpose: Returns field Ranking
    SetRanking (me: mutable; Ranking: Integer);
	---Purpose: Set field Ranking

    RankingRationale (me) returns HAsciiString from TCollection;
	---Purpose: Returns field RankingRationale
    SetRankingRationale (me: mutable; RankingRationale: HAsciiString from TCollection);
	---Purpose: Set field RankingRationale

    Quantity (me) returns MeasureWithUnit from StepBasic;
	---Purpose: Returns field Quantity
    SetQuantity (me: mutable; Quantity: MeasureWithUnit from StepBasic);
	---Purpose: Set field Quantity

fields
    theRanking: Integer;
    theRankingRationale: HAsciiString from TCollection;
    theQuantity: MeasureWithUnit from StepBasic;

end MakeFromUsageOption;
