-- File:	StepToTopoDS_TranslateVertex.cdl
-- Created:	Fri Dec 16 14:48:28 1994
-- Author:	Frederic MAUPAS
--		<fma@stylox>
---Copyright:	 Matra Datavision 1994

class TranslateVertex from StepToTopoDS
    inherits Root from StepToTopoDS
    
    ---Purpose:
    --         

uses

    Vertex               from StepShape,
    TranslateVertexError from StepToTopoDS,
    Tool                 from StepToTopoDS,
    Shape                from TopoDS,
    NMTool               from StepToTopoDS

raises NotDone from StdFail

is

    Create returns TranslateVertex;
    
    Create (V      : Vertex        from StepShape;
            T      : in out Tool   from StepToTopoDS;
            NMTool : in out NMTool from StepToTopoDS)
    	returns TranslateVertex;
	    
    Init (me     : in out;
          V      : Vertex        from StepShape;
          T      : in out Tool   from StepToTopoDS;
          NMTool : in out NMTool from StepToTopoDS);

    Value (me) returns Shape from TopoDS
    	raises NotDone
	is static;
	---C++: return const &

    Error (me) returns TranslateVertexError from StepToTopoDS;
    
fields

    myError  : TranslateVertexError from StepToTopoDS;
    
    myResult : Shape                from TopoDS;
    
end TranslateVertex;
