-- File:	StepToGeom_MakeVectorWithMagnitude.cdl
-- Created:	Mon Jun 14 15:10:06 1993
-- Author:	Martine LANGLOIS
---Copyright:	 Matra Datavision 1993

class MakeVectorWithMagnitude from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          Vector from StepGeom which describes a VectorWithMagnitude 
    --          from Prostep and VectorWithMagnitude from Geom.

uses 
     VectorWithMagnitude from Geom,
     Vector from StepGeom

is 

    Convert ( myclass; SV : Vector from StepGeom;
                       CV : out VectorWithMagnitude from Geom )
    returns Boolean from Standard;

end MakeVectorWithMagnitude;
