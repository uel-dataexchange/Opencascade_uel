-- File:	GeomToStep_MakeBSplineCurveWithKnotsAndRationalBSplineCurve.cdl
-- Created:	Mon Jun 14 15:22:02 1993
-- Author:	Martine LANGLOIS
--		<mla@mastox>
---Copyright:	 Matra Datavision 1993

class MakeBSplineCurveWithKnotsAndRationalBSplineCurve from GeomToStep inherits
    Root from GeomToStep

    ---Purpose: This class implements the mapping between classes
    --          BSplineCurve from Geom, Geom2d and the class
    --          BSplineCurveWithKnotsAndRationalBSplineCurve from StepGeom
    --          which describes a rational_bspline_curve_with_knots from
    --          Prostep
  
uses

     BSplineCurve from Geom,
     BSplineCurve from Geom2d,
     BSplineCurveWithKnotsAndRationalBSplineCurve from StepGeom
     
raises

     NotDone from StdFail
     
is 

Create ( Bsplin : BSplineCurve from Geom ) returns
    MakeBSplineCurveWithKnotsAndRationalBSplineCurve;

Create ( Bsplin : BSplineCurve from Geom2d ) returns
    MakeBSplineCurveWithKnotsAndRationalBSplineCurve;
Value (me) returns
    BSplineCurveWithKnotsAndRationalBSplineCurve from StepGeom
    raises NotDone
    is static;
    ---C++: return const&
    
fields

    theBSplineCurveWithKnotsAndRationalBSplineCurve :
    	BSplineCurveWithKnotsAndRationalBSplineCurve from StepGeom;
    	-- The solution from StepGeom
    	
end MakeBSplineCurveWithKnotsAndRationalBSplineCurve;
