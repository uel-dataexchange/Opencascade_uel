-- File:	GeomToStep_MakeSurfaceOfLinearExtrusion.cdl
-- Created:	Mon Jun 14 16:16:49 1993
-- Author:	Martine LANGLOIS
--		<mla@mastox>
---Copyright:	 Matra Datavision 1993

class MakeSurfaceOfLinearExtrusion from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between class
    --          SurfaceOfLinearExtrusion from Geom and the class
    --          SurfaceOfLinearExtrusion from StepGeom which describes a
    --          surface_of_linear_extrusion from Prostep
  
uses SurfaceOfLinearExtrusion from Geom,
     SurfaceOfLinearExtrusion from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( CSurf : SurfaceOfLinearExtrusion from Geom ) returns
    MakeSurfaceOfLinearExtrusion;

Value (me) returns SurfaceOfLinearExtrusion from StepGeom
    raises NotDone
    is static;
    ---C++: return const&

fields

    theSurfaceOfLinearExtrusion : SurfaceOfLinearExtrusion from StepGeom;
    	-- The solution from StepGeom
    	
end MakeSurfaceOfLinearExtrusion;


