-- File:	IGESAppli_ToolPinNumber.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolPinNumber  from IGESAppli

    ---Purpose : Tool to work on a PinNumber. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses PinNumber from IGESAppli,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolPinNumber;
    ---Purpose : Returns a ToolPinNumber, ready to work


    ReadOwnParams (me; ent : mutable PinNumber;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : PinNumber;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : PinNumber;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a PinNumber <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable PinNumber) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a PinNumber
    --           (Level cleared in D.E. if Subordinate != 0)

    DirChecker (me; ent : PinNumber) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : PinNumber;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : PinNumber; entto : mutable PinNumber;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : PinNumber;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolPinNumber;
