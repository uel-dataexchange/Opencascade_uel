-- File:	TopOpeBRepBuild_ShellToSolid.cdl
-- Created:	Thu Oct  2 15:17:26 1997
-- Author:	Xuan Trang PHAM PHU
--		<xpu@poulopox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


class ShellToSolid from TopOpeBRepBuild

---Purpose: 
-- This class builds solids from a set of shells SSh and a solid F. 

uses

    Shell from TopoDS,
    Solid from TopoDS,
    ListOfShape from TopTools

is

    Create returns ShellToSolid;
     
    Init(me : in out)
    is static;
    
    AddShell(me : in out; Sh : Shell from TopoDS)
    is  static;
     	
    MakeSolids(me : in out; 
    	       So : Solid from TopoDS;
    	       LSo : in out ListOfShape from TopTools)
    is static;

fields 

    myLSh : ListOfShape from TopTools;
    
end ShellToSolid;
