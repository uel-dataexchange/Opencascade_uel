-- File:	IGESGraph_ToolLineFontPredefined.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolLineFontPredefined  from IGESGraph

    ---Purpose : Tool to work on a LineFontPredefined. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses LineFontPredefined from IGESGraph,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolLineFontPredefined;
    ---Purpose : Returns a ToolLineFontPredefined, ready to work


    ReadOwnParams (me; ent : mutable LineFontPredefined;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : LineFontPredefined;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : LineFontPredefined;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a LineFontPredefined <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable LineFontPredefined) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a LineFontPredefined
    --           (NbPropertyValues forced to 1)

    DirChecker (me; ent : LineFontPredefined) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : LineFontPredefined;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : LineFontPredefined; entto : mutable LineFontPredefined;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : LineFontPredefined;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolLineFontPredefined;
