-- File:	RWStepShape_RWAngularLocation.cdl
-- Created:	Tue Apr 18 16:42:57 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWAngularLocation from RWStepShape

    ---Purpose: Read & Write tool for AngularLocation

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    AngularLocation from StepShape

is
    Create returns RWAngularLocation from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : AngularLocation from StepShape);
	---Purpose: Reads AngularLocation

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: AngularLocation from StepShape);
	---Purpose: Writes AngularLocation

    Share (me; ent : AngularLocation from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWAngularLocation;
