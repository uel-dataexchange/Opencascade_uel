-- File:	RWStepDimTol_RWLineProfileTolerance.cdl
-- Created:	Wed Jun  4 13:34:34 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWLineProfileTolerance from RWStepDimTol

    ---Purpose: Read & Write tool for LineProfileTolerance

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    LineProfileTolerance from StepDimTol

is
    Create returns RWLineProfileTolerance from RWStepDimTol;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : LineProfileTolerance from StepDimTol);
	---Purpose: Reads LineProfileTolerance

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: LineProfileTolerance from StepDimTol);
	---Purpose: Writes LineProfileTolerance

    Share (me; ent : LineProfileTolerance from StepDimTol;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWLineProfileTolerance;
