-- File:	TDF_ChildIDIterator.cdl
--      	-----------------------
-- Author:	DAUTRY Philippe
--		<fid@fox.paris1.matra-dtv.fr>
---Copyright:	 MATRA DATAVISION 1997

---Version:	0.0
---History:	Version	Date		Purpose
--		0.0	Nov 20 1997	Creation

class ChildIDIterator from TDF 

	---Purpose: Iterates on the children of a label, to find
	--          attributes having ID as Attribute ID.
	--          
	--          Level option works as TDF_ChildIterator.

uses

    Attribute     from TDF,
    Label         from TDF,
    LabelNodePtr  from TDF,
    ChildIterator from TDF
    
is

    Create
    	returns ChildIDIterator from TDF;
    	---Purpose: Creates an empty iterator.
    
    Create(aLabel    : Label from TDF;
    	   anID      : GUID from Standard;
    	   allLevels : Boolean from Standard = Standard_False)
    	returns ChildIDIterator from TDF;
    	---Purpose: Iterates on the children of the given label. If
    	--          <allLevels> option is set to true, it explores not
    	--          only the first, but all the sub label levels.
    
    Initialize(me : in out;
    	       aLabel    : Label from TDF;
    	       anID      : GUID from Standard;
    	       allLevels : Boolean from Standard = Standard_False);
    	---Purpose: Initializes the iteration on the children of the
    	--          given label. If <allLevels> option is set to true,
    	--          it explores not only the first, but all the sub
    	--          label levels.
    
    More(me) returns Boolean;
	---Purpose: Returns True if there is a current Item in the
	--          iteration.
	--          
	---C++: inline

    Next(me : in out);
    	---Purpose: Move to the next Item 
    
    NextBrother(me : in out);
    	---Purpose: Move to the next Brother. If there is none, go up
    	--          etc. This method is interesting only with
    	--          "allLevels" behavior, because it avoids to explore
    	--          the current label children.
    
    Value(me) returns Attribute from TDF;
	---Purpose: Returns the current item; a null handle if there is none.
	--          
	---C++: inline

fields

    myID  : GUID from Standard;
    myItr : ChildIterator  from TDF;
    myAtt : Attribute from TDF;

end ChildIDIterator;
