-- File:	StepBasic_Action.cdl
-- Created:	Fri Nov 26 16:26:28 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class Action from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity Action

uses
    HAsciiString from TCollection,
    ActionMethod from StepBasic

is
    Create returns Action from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       hasDescription: Boolean;
                       aDescription: HAsciiString from TCollection;
                       aChosenMethod: ActionMethod from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description
    HasDescription (me) returns Boolean;
	---Purpose: Returns True if optional field Description is defined

    ChosenMethod (me) returns ActionMethod from StepBasic;
	---Purpose: Returns field ChosenMethod
    SetChosenMethod (me: mutable; ChosenMethod: ActionMethod from StepBasic);
	---Purpose: Set field ChosenMethod

fields
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection; -- optional
    theChosenMethod: ActionMethod from StepBasic;
    defDescription: Boolean; -- flag "is Description defined"

end Action;
