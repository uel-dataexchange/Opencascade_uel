-- File:	RWStepBasic_RWRoleAssociation.cdl
-- Created:	Wed May 10 15:09:08 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWRoleAssociation from RWStepBasic

    ---Purpose: Read & Write tool for RoleAssociation

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    RoleAssociation from StepBasic

is
    Create returns RWRoleAssociation from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : RoleAssociation from StepBasic);
	---Purpose: Reads RoleAssociation

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: RoleAssociation from StepBasic);
	---Purpose: Writes RoleAssociation

    Share (me; ent : RoleAssociation from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWRoleAssociation;
