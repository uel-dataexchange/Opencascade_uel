-- File:	MakeHyperbola.cdl
-- Created:	Mon Sep 28 11:49:29 1992
-- Author:	Remi GILET
--		<reg@sdsun2>
---Copyright:	 Matra Datavision 1992

class MakeHyperbola from GC inherits Root from GC

    ---Purpose :This class implements construction algorithms for a hyperbola in
    -- 3D space. The result is a Geom_Hyperbola hyperbola.
    -- A MakeHyperbola object provides a framework for:
    -- -   defining the construction of the hyperbola,
    -- -   implementing the construction algorithm, and
    -- -   consulting the results. In particular, the Value
    --   function returns the constructed hyperbola.
    --  To define the main branch of an hyperbola.
    --  The parameterization range is ]-infinite,+infinite[
    --  It is possible to get the other branch and the two conjugate
    --  branches of the main branch.
    --
    --                         ^YAxis                
    --                         |                   
    --                  FirstConjugateBranch     
    --                         |        
    --        Other            |                Main
    --   --------------------- C ------------------------------>XAxis
    --        Branch           |                Branch
    --                         |         
    --                   SecondConjugateBranch
    --                         |         
    --
    --  The major radius is the distance between the Location point
    --  of the hyperbola C and the apex of the Main Branch (or the
    --  Other branch). The major axis is the XAxis.
    --  The minor radius is the distance between the Location point
    --  of the hyperbola C and the apex of the First (or Second)
    --  Conjugate branch. The minor axis is the YAxis.
    --  The major radius can be lower than the minor radius.

uses Pnt       from gp,
     Hypr      from gp,
     Ax2       from gp,
     Hyperbola from Geom

raises NotDone from StdFail

is

Create (H : Hypr from gp)   returns MakeHyperbola;
    --- Purpose :
    --  Creates  an Hyperbola from a non persistent hyperbola  from package gp by conversion.

Create (A2 : Ax2                        from gp      ; 
    	MajorRadius, MinorRadius : Real from Standard) returns MakeHyperbola;
    --- Purpose : Constructs a hyperbola centered on the origin of the coordinate system
    -- A2, with major and minor radii MajorRadius and MinorRadius, where:
    --   the plane of the hyperbola is defined by the "X Axis" and "Y Axis" of A2,
    --   -   its major axis is the "X Axis" of A2.

Create(S1,S2  : Pnt from gp;
       Center : Pnt from gp) returns MakeHyperbola;
    ---Purpose: Constructs a hyperbola centered on the point Center, where
    --   -   the plane of the hyperbola is defined by Center, S1 and S2,
    --   -   its major axis is defined by Center and S1,
    --   -   its major radius is the distance between Center and S1, and
    --   -   its minor radius is the distance between S2 and the major axis;
		
Value(me) returns Hyperbola from Geom
    raises NotDone
    is static;
    ---Purpose: Returns the constructed hyperbola.
    -- Exceptions StdFail_NotDone if no hyperbola is constructed.
    ---C++: return const&

Operator(me) returns Hyperbola from Geom
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator Handle_Geom_Hyperbola() const;"

fields

    TheHyperbola : Hyperbola from Geom;
    --The solution from Geom.
    
end MakeHyperbola;
