-- File:	StepRepr_Extension.cdl
-- Created:	Tue Apr 24 13:47:10 2001
-- Author:	Christian CAILLET
--		<cky@photox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 2001

class Extension  from StepRepr    inherits DerivedShapeAspect  from StepRepr

    ---Purpose : Added for Dimensional Tolerances

uses
    Integer

is

    Create returns mutable Extension;

end Extension;
