-- File:	StepRepr_ProductDefinitionUsage.cdl
-- Created:	Mon Jul  3 19:47:51 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class ProductDefinitionUsage from StepRepr
inherits ProductDefinitionRelationship from StepBasic

    ---Purpose: Representation of STEP entity ProductDefinitionUsage

uses
    HAsciiString from TCollection,
    ProductDefinition from StepBasic

is
    Create returns ProductDefinitionUsage from StepRepr;
	---Purpose: Empty constructor

end ProductDefinitionUsage;
