-- File:	StepAP214_AppliedExternalIdentificationAssignment.cdl
-- Created:	Wed May 10 15:09:06 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class AppliedExternalIdentificationAssignment from StepAP214
inherits ExternalIdentificationAssignment from StepBasic

    ---Purpose: Representation of STEP entity AppliedExternalIdentificationAssignment

uses
    HAsciiString from TCollection,
    IdentificationRole from StepBasic,
    ExternalSource from StepBasic,
    HArray1OfExternalIdentificationItem from StepAP214

is
    Create returns AppliedExternalIdentificationAssignment from StepAP214;
	---Purpose: Empty constructor

    Init (me: mutable; aIdentificationAssignment_AssignedId: HAsciiString from TCollection;
                       aIdentificationAssignment_Role: IdentificationRole from StepBasic;
                       aExternalIdentificationAssignment_Source: ExternalSource from StepBasic;
                       aItems: HArray1OfExternalIdentificationItem from StepAP214);
	---Purpose: Initialize all fields (own and inherited)

    Items (me) returns HArray1OfExternalIdentificationItem from StepAP214;
	---Purpose: Returns field Items
    SetItems (me: mutable; Items: HArray1OfExternalIdentificationItem from StepAP214);
	---Purpose: Set field Items

fields
    theItems: HArray1OfExternalIdentificationItem from StepAP214;

end AppliedExternalIdentificationAssignment;
