-- File:	IGESGeom_ToolCurveOnSurface.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolCurveOnSurface  from IGESGeom

    ---Purpose : Tool to work on a CurveOnSurface. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses CurveOnSurface from IGESGeom,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolCurveOnSurface;
    ---Purpose : Returns a ToolCurveOnSurface, ready to work


    ReadOwnParams (me; ent : mutable CurveOnSurface;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : CurveOnSurface;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : CurveOnSurface;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a CurveOnSurface <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable CurveOnSurface) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a CurveOnSurface
    --           (its CurveUV must have UseFlag at 5)

    DirChecker (me; ent : CurveOnSurface) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : CurveOnSurface;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : CurveOnSurface; entto : mutable CurveOnSurface;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : CurveOnSurface;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolCurveOnSurface;
