-- File:	Geom2dToIGES.cdl
-- Created:	Thu Nov 17 13:55:58 1994
-- Author:	Marie Jose MARTZ
--		<mjm@minox>
---Copyright:	 Matra Datavision 1994

package Geom2dToIGES

--- Purpose: Creation des entites geometriques de IGES
--           a partir des entites de Geom2d.

uses Interface, IGESData, IGESBasic, IGESConvGeom, IGESGeom, IGESSolid, IGESToBRep,
     gp, Geom, Geom2d, GeomLProp, TColStd, TopoDS, TopTools,
     Transfer, TransferBRep, BRep, TCollection, ElCLib

is

-- classes du package

    class Geom2dCurve;
    class Geom2dEntity;
    class Geom2dPoint;    
    class Geom2dVector;


end Geom2dToIGES;
