-- File:        PresentationStyleByContext.cdl
-- Created:     Fri Dec  1 11:11:25 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class PresentationStyleByContext from StepVisual 

inherits PresentationStyleAssignment from StepVisual 

uses

	StyleContextSelect from StepVisual, 
	HArray1OfPresentationStyleSelect from StepVisual
is

	Create returns mutable PresentationStyleByContext;
	---Purpose: Returns a PresentationStyleByContext


	Init (me : mutable;
	      aStyles : mutable HArray1OfPresentationStyleSelect from StepVisual) is redefined;

	Init (me : mutable;
	      aStyles : mutable HArray1OfPresentationStyleSelect from StepVisual;
	      aStyleContext : StyleContextSelect from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetStyleContext(me : mutable; aStyleContext : StyleContextSelect);
	StyleContext (me) returns StyleContextSelect;

fields

	styleContext : StyleContextSelect from StepVisual; -- a SelectType

end PresentationStyleByContext;
