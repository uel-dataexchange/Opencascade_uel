-- File:        CsgPrimitive.cdl
-- Created:     Fri Dec  1 11:11:10 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class CsgPrimitive from StepShape inherits SelectType from StepData

	-- <CsgPrimitive> is an EXPRESS Select Type construct translation.
	-- it gathers : Sphere, Block, RightAngularWedge, Torus, RightCircularCone, RightCircularCylinder

uses

	Sphere,
	Block,
	RightAngularWedge,
	Torus,
	RightCircularCone,
	RightCircularCylinder
is

	Create returns CsgPrimitive;
	---Purpose : Returns a CsgPrimitive SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a CsgPrimitive Kind Entity that is :
	--        1 -> Sphere
	--        2 -> Block
	--        3 -> RightAngularWedge
	--        4 -> Torus
	--        5 -> RightCircularCone
	--        6 -> RightCircularCylinder
	--        0 else

	Sphere (me) returns any Sphere;
	---Purpose : returns Value as a Sphere (Null if another type)

	Block (me) returns any Block;
	---Purpose : returns Value as a Block (Null if another type)

	RightAngularWedge (me) returns any RightAngularWedge;
	---Purpose : returns Value as a RightAngularWedge (Null if another type)

	Torus (me) returns any Torus;
	---Purpose : returns Value as a Torus (Null if another type)

	RightCircularCone (me) returns any RightCircularCone;
	---Purpose : returns Value as a RightCircularCone (Null if another type)

	RightCircularCylinder (me) returns any RightCircularCylinder;
	---Purpose : returns Value as a RightCircularCylinder (Null if another type)


end CsgPrimitive;

