-- File:	PCollection_Hash.cdl
-- Created:	Mon Apr 22 16:26:20 1991
-- Author:	jean pierre TIRAULT
--		<jpt@topsn1>
---Copyright:	 Matra Datavision 1991


generic class Hash from PCollection (key as Storable) inherits Storable
    is
    
    
    
    Create returns Hash;
    ---Purpose : Empty constructor.



    HashCode (me; MyKey : key ; Upper : Integer) 
             returns Integer is virtual;
    ---Level: Public
    ---Purpose: Returns a hashcod value of key bounded by Upper.



    Compare (me; One , Two : key) returns Boolean is virtual;    
    ---Level: Public
    ---Purpose : Compare two keys and returns a boolean value

end;

