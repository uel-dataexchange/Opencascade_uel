-- File:	RWStepAP214_RWAppliedExternalIdentificationAssignment.cdl
-- Created:	Wed May 10 15:09:06 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWAppliedExternalIdentificationAssignment from RWStepAP214

    ---Purpose: Read & Write tool for AppliedExternalIdentificationAssignment

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    AppliedExternalIdentificationAssignment from StepAP214

is
    Create returns RWAppliedExternalIdentificationAssignment from RWStepAP214;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : AppliedExternalIdentificationAssignment from StepAP214);
	---Purpose: Reads AppliedExternalIdentificationAssignment

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: AppliedExternalIdentificationAssignment from StepAP214);
	---Purpose: Writes AppliedExternalIdentificationAssignment

    Share (me; ent : AppliedExternalIdentificationAssignment from StepAP214;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWAppliedExternalIdentificationAssignment;
