-- File:	RWStepRepr_RWQuantifiedAssemblyComponentUsage.cdl
-- Created:	Mon Jul  3 20:13:37 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWQuantifiedAssemblyComponentUsage from RWStepRepr

    ---Purpose: Read & Write tool for QuantifiedAssemblyComponentUsage

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    QuantifiedAssemblyComponentUsage from StepRepr

is
    Create returns RWQuantifiedAssemblyComponentUsage from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : QuantifiedAssemblyComponentUsage from StepRepr);
	---Purpose: Reads QuantifiedAssemblyComponentUsage

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: QuantifiedAssemblyComponentUsage from StepRepr);
	---Purpose: Writes QuantifiedAssemblyComponentUsage

    Share (me; ent : QuantifiedAssemblyComponentUsage from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWQuantifiedAssemblyComponentUsage;
