-- File:	HLRTest_Projector.cdl
-- Created:	Wed Apr  5 16:30:59 1995
-- Author:	Christophe MARION
--		<cma@ecolox>
---Copyright:	 Matra Datavision 1995

class Projector from HLRTest inherits Drawable3D from Draw
	---Purpose: 

uses
    OStream,
    Display     from Draw,
    Interpretor from Draw,
    Projector   from HLRAlgo

is
    Create(P : Projector from HLRAlgo)
    returns mutable Projector from HLRTest; 
    
    Projector(me) returns Projector from HLRAlgo;
	---C++: return const &
	---C++: inline

    DrawOn(me; dis : in out Display from Draw);
	---Purpose: Does nothhing,
    
    Copy(me) returns mutable Drawable3D from Draw
	---Purpose: For variable copy.
    is redefined;
	
    Dump(me; S : in out OStream)
	---Purpose: For variable dump.
    is redefined;

    Whatis(me; I : in out Interpretor from Draw)
	---Purpose: For variable whatis command. Set  as a result  the
	--          type of the variable.
    is redefined;

fields
    myProjector : Projector from HLRAlgo;

end Projector;
