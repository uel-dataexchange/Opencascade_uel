-- File:        ReversibleTopologyItem.cdl
-- Created:     Fri Dec  1 11:11:11 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class ReversibleTopologyItem from StepShape inherits SelectType from StepData

	-- <ReversibleTopologyItem> is an EXPRESS Select Type construct translation.
	-- it gathers : Edge, Path, Face, FaceBound, ClosedShell, OpenShell

uses

	Edge,
	Path,
	Face,
	FaceBound,
	ClosedShell,
	OpenShell
is

	Create returns ReversibleTopologyItem;
	---Purpose : Returns a ReversibleTopologyItem SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a ReversibleTopologyItem Kind Entity that is :
	--        1 -> Edge
	--        2 -> Path
	--        3 -> Face
	--        4 -> FaceBound
	--        5 -> ClosedShell
	--        6 -> OpenShell
	--        0 else

	Edge (me) returns any Edge;
	---Purpose : returns Value as a Edge (Null if another type)

	Path (me) returns any Path;
	---Purpose : returns Value as a Path (Null if another type)

	Face (me) returns any Face;
	---Purpose : returns Value as a Face (Null if another type)

	FaceBound (me) returns any FaceBound;
	---Purpose : returns Value as a FaceBound (Null if another type)

	ClosedShell (me) returns any ClosedShell;
	---Purpose : returns Value as a ClosedShell (Null if another type)

	OpenShell (me) returns any OpenShell;
	---Purpose : returns Value as a OpenShell (Null if another type)


end ReversibleTopologyItem;

