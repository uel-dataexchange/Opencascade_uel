-- File:        FacetedBrepShapeRepresentation.cdl
-- Created:     Mon Dec  4 12:02:27 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWFacetedBrepShapeRepresentation from RWStepShape

	---Purpose : Read & Write Module for FacetedBrepShapeRepresentation

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     FacetedBrepShapeRepresentation from StepShape,
     EntityIterator from Interface

is

	Create returns RWFacetedBrepShapeRepresentation;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable FacetedBrepShapeRepresentation from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : FacetedBrepShapeRepresentation from StepShape);

	Share(me; ent : FacetedBrepShapeRepresentation from StepShape; iter : in out EntityIterator);

end RWFacetedBrepShapeRepresentation;
