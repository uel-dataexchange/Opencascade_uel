-- File:	RWStepRepr_RWConfigurationDesign.cdl
-- Created:	Fri Nov 26 16:26:36 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWConfigurationDesign from RWStepRepr

    ---Purpose: Read & Write tool for ConfigurationDesign

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ConfigurationDesign from StepRepr

is
    Create returns RWConfigurationDesign from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ConfigurationDesign from StepRepr);
	---Purpose: Reads ConfigurationDesign

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ConfigurationDesign from StepRepr);
	---Purpose: Writes ConfigurationDesign

    Share (me; ent : ConfigurationDesign from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWConfigurationDesign;
