-- File:	GeomFill_Profiler.cdl
-- Created:	Thu Feb 17 10:44:36 1994
-- Author:	Bruno DUMORTIER
--		<dub@fuegox>
---Copyright:	 Matra Datavision 1994




class Profiler from GeomFill

	---Purpose: Evaluation of the common BSplineProfile of a group
	--          of curves  from Geom. All the curves will have the
	--          same  degree,  the same knot-vector, so  the  same
	--          number of poles.


uses
    Array1OfReal    from TColStd,
    Array1OfInteger from TColStd,
    Array1OfPnt     from TColgp,
    Curve           from Geom,
    SequenceOfCurve from TColGeom


raises
    NotDone     from StdFail,
    DomainError from Standard

is
    Create returns Profiler from GeomFill;
    
    Delete(me:out) is virtual;
    ---C++: alias "Standard_EXPORT virtual ~GeomFill_Profiler(){Delete() ; }"
    
    AddCurve( me    : in out;
              Curve : in Curve from Geom)
    is static;
    
    Perform(me   : in out ;
            PTol : in Real from Standard)
	---Purpose: Converts all curves to BSplineCurves.
	--          Set them to the common profile.
	--          <PTol> is used to compare 2 knots.
    is virtual;
    
    Degree(me) returns Integer from Standard
    raises 
    	NotDone from StdFail
	---Purpose: Raises if not yet perform
    is static;
    
    IsPeriodic(me) returns Boolean from Standard
	---C++: inline
    is static;
    
    NbPoles(me) returns Integer from Standard
    raises 
    	NotDone from StdFail
	---Purpose: Raises if not yet perform
    is static;
    
    Poles(me; Index : in     Integer     from Standard;
    	      Poles : in out Array1OfPnt from TColgp)
    	---Purpose: returns in <Poles> the  poles  of the BSplineCurve
    	--          from index <Index> adjusting to the current profile.
    raises 
    	NotDone     from StdFail,
	---Purpose: Raises if not yet perform
    	DomainError from Standard
	---Purpose: Raises if <Index> not in the range [1,NbCurves]
	--          if  the  length  of  <Poles>  is  not  equal  to
	--          NbPoles().
    is static;
    
    Weights(me; Index   : in     Integer      from Standard;
    	        Weights : in out Array1OfReal from TColStd)
    	---Purpose: returns in <Weights> the weights of the BSplineCurve
    	--          from index <Index> adjusting to the current profile.
    raises 
    	NotDone from StdFail,
	---Purpose: Raises if not yet perform
    	DomainError from Standard
	---Purpose: Raises if <Index> not in the range [1,NbCurves] or
	--          if  the  length  of  <Weights>  is  not  equal  to
	--          NbPoles().
    is static;
    
    NbKnots(me) returns Integer from Standard
    raises 
    	NotDone from StdFail
	---Purpose: Raises if not yet perform
    is static;
    
    KnotsAndMults(me;
                  Knots : in out Array1OfReal    from TColStd;
		  Mults : in out Array1OfInteger from TColStd)
    raises 
    	NotDone from StdFail,
	---Purpose: Raises if not yet perform
    	DomainError from Standard
	---Purpose: Raises if  the lengthes of <Knots> and <Mults> are
	--          not equal to NbKnots().
    is static;
    
    Curve(me; Index : Integer from Standard) 
    returns Curve from Geom
    	---C++: return const&
    	---C++: inline
    is static;
    
    
fields
    mySequence   : SequenceOfCurve from TColGeom is protected;
    myIsDone     : Boolean         from Standard is protected;
    myIsPeriodic : Boolean         from Standard is protected;

end Profiler;
