-- File:        OrientedOpenShell.cdl
-- Created:     Fri Dec  1 11:11:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class OrientedOpenShell from StepShape 

inherits OpenShell from StepShape 

uses

	Boolean from Standard, 
	HArray1OfFace from StepShape, 
	Face from StepShape, 
	HAsciiString from TCollection
is

	Create returns mutable OrientedOpenShell;
	---Purpose: Returns a OrientedOpenShell


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aCfsFaces : mutable HArray1OfFace from StepShape) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aOpenShellElement : mutable OpenShell from StepShape;
	      aOrientation : Boolean from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetOpenShellElement(me : mutable; aOpenShellElement : mutable OpenShell);
	OpenShellElement (me) returns mutable OpenShell;
	SetOrientation(me : mutable; aOrientation : Boolean);
	Orientation (me) returns Boolean;
	SetCfsFaces(me : mutable; aCfsFaces : mutable HArray1OfFace) is redefined;
	CfsFaces (me) returns mutable HArray1OfFace is redefined;
	CfsFacesValue (me; num : Integer) returns mutable Face is redefined;
	NbCfsFaces (me) returns Integer is redefined;

fields

	openShellElement : OpenShell from StepShape;
	orientation : Boolean from Standard;

 -- 
 -- NB : field <cfs_faces> inherited from classe <connected_face_set> is redeclared.
 --      it shall appears in a physical file as a *.
 --

end OrientedOpenShell;
