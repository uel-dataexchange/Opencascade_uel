-- File:	BinDrivers.cdl
-- Created:	Tue Oct 29 11:30:48 2002
-- Author:	Michael SAZONOV
--		<msv@novgorox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2002


package BinDrivers

uses
    Standard,
    TDF,
    TCollection,
    TColStd,
    CDM,
    PCDM,
    Storage,
    BinObjMgt,
    BinMDF,
    BinLDrivers

is

    class DocumentStorageDriver;
    class DocumentRetrievalDriver;

    Factory (theGUID : GUID from Standard) returns Transient from Standard;

    AttributeDrivers (MsgDrv : MessageDriver from CDM)
    	returns ADriverTable from BinMDF;
    	---Purpose: Creates the table of drivers of types supported

    StorageVersion returns AsciiString from TCollection;
        ---Purpose: returns "1"
    
end BinDrivers;
