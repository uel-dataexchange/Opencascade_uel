-- File:	StepToTopoDS_GeometricTool.cdl
-- Created:	Thu Jan  5 15:56:59 1995
-- Author:	Frederic MAUPAS
--		<fma@stylox>
---Copyright:	 Matra Datavision 1995

class GeometricTool from StepToTopoDS

  ---Purpose: This class contains some algorithmic services 
  --          specific to the mapping STEP to CAS.CADE              

uses

    Tool         from StepToTopoDS,
    SurfaceCurve from StepGeom,
    Surface      from StepGeom,
    Pcurve       from StepGeom,
    EdgeLoop     from StepShape,    
    Edge         from StepShape,    
    Curve        from Geom2d,
    Line         from Geom2d,
    Curve        from Geom,
    Surface      from Geom,
    Pnt2d        from gp,
    Pnt          from gp,
    Face         from TopoDS,
    Wire         from TopoDS,
    Edge         from TopoDS,
    Vertex       from TopoDS
    
is

    PCurve(myclass;
 	      SC : SurfaceCurve from StepGeom;
    	      S  : Surface      from StepGeom;
	      PC : out Pcurve   from StepGeom;
	      last : Integer = 0)
    	returns Integer;

    IsSeamCurve(myclass;
    	    	SC : SurfaceCurve from StepGeom;
    	      	S  : Surface      from StepGeom;
		E  : Edge         from StepShape;
    	    	EL : EdgeLoop     from StepShape)
    	returns Boolean;

		
    IsLikeSeam(myclass;
    	       SC : SurfaceCurve from StepGeom;
       	       S  : Surface      from StepGeom;
	       E  : Edge         from StepShape;
    	       EL : EdgeLoop     from StepShape)
    	returns Boolean;


    UpdateParam3d(myclass; C  : Curve from Geom;
    	    	  w1, w2 : in out Real from Standard;
		  preci  : Real)
    	returns Boolean;
			 
end GeometricTool from StepToTopoDS;
