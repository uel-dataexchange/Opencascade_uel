-- File:        QualifiedRepresentationItem.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWQualifiedRepresentationItem from RWStepShape

	---Purpose : Read & Write Module for QualifiedRepresentationItem

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     QualifiedRepresentationItem from StepShape,
     EntityIterator from Interface

is

	Create returns RWQualifiedRepresentationItem;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable QualifiedRepresentationItem from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : QualifiedRepresentationItem from StepShape);

	Share(me; ent : QualifiedRepresentationItem from StepShape; iter : in out EntityIterator);

end RWQualifiedRepresentationItem;
