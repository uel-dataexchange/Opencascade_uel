-- File:        TrimmedCurve.cdl
-- Created:     Mon Dec  4 12:02:32 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWTrimmedCurve from RWStepGeom

	---Purpose : Read & Write Module for TrimmedCurve

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     TrimmedCurve from StepGeom,
     EntityIterator from Interface

is

	Create returns RWTrimmedCurve;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable TrimmedCurve from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : TrimmedCurve from StepGeom);

	Share(me; ent : TrimmedCurve from StepGeom; iter : in out EntityIterator);

end RWTrimmedCurve;
