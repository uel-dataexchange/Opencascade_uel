-- File:	IGESDimen_ToolOrdinateDimension.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolOrdinateDimension  from IGESDimen

    ---Purpose : Tool to work on a OrdinateDimension. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses OrdinateDimension from IGESDimen,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolOrdinateDimension;
    ---Purpose : Returns a ToolOrdinateDimension, ready to work


    ReadOwnParams (me; ent : mutable OrdinateDimension;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : OrdinateDimension;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : OrdinateDimension;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a OrdinateDimension <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : OrdinateDimension) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : OrdinateDimension;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : OrdinateDimension; entto : mutable OrdinateDimension;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : OrdinateDimension;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolOrdinateDimension;
