-- File:	IGESDimen_ToolDiameterDimension.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolDiameterDimension  from IGESDimen

    ---Purpose : Tool to work on a DiameterDimension. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses DiameterDimension from IGESDimen,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolDiameterDimension;
    ---Purpose : Returns a ToolDiameterDimension, ready to work


    ReadOwnParams (me; ent : mutable DiameterDimension;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : DiameterDimension;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : DiameterDimension;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a DiameterDimension <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : DiameterDimension) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : DiameterDimension;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : DiameterDimension; entto : mutable DiameterDimension;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : DiameterDimension;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolDiameterDimension;
