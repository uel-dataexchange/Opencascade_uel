-- File:        PlaneAngleUnit.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPlaneAngleUnit from RWStepBasic

	---Purpose : Read & Write Module for PlaneAngleUnit

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PlaneAngleUnit from StepBasic,
     EntityIterator from Interface

is

	Create returns RWPlaneAngleUnit;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PlaneAngleUnit from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : PlaneAngleUnit from StepBasic);

	Share(me; ent : PlaneAngleUnit from StepBasic; iter : in out EntityIterator);

end RWPlaneAngleUnit;
