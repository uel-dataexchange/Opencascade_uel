-- File:        BooleanResult.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWBooleanResult from RWStepShape

	---Purpose : Read & Write Module for BooleanResult

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     BooleanResult from StepShape,
     EntityIterator from Interface

is

	Create returns RWBooleanResult;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable BooleanResult from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : BooleanResult from StepShape);

	Share(me; ent : BooleanResult from StepShape; iter : in out EntityIterator);

end RWBooleanResult;
