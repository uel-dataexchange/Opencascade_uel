-- File:	AppCont_TheLineTool.cdl
-- Created:	Thu Apr 22 12:02:11 1993
-- Author:	Laurent PAINNOT
--		<lpa@phobox>
---Copyright:	 Matra Datavision 1993


deferred generic class TheLineTool from AppCont(MLine as any)

    ---Purpose: Template for desribing a continuous MultiLine.
    --          The Vectors returned by the methods Tangency are
    --          the derivative values.

uses
     Pnt           from gp,
     Pnt2d         from gp,
     Vec           from gp,
     Vec2d         from gp,
     Array1OfPnt   from TColgp,
     Array1OfPnt2d from TColgp,
     Array1OfVec   from TColgp,
     Array1OfVec2d from TColgp

is
    
    FirstParameter(myclass; ML: MLine) returns Real;
    	---Purpose: returns the first parameter of the Line.

    LastParameter(myclass; ML: MLine) returns Real;
    	---Purpose: returns the last parameter of the Line.

    NbP2d(myclass; ML: MLine) returns Integer;
    	---Purpose: Returns the number of 2d points of a MLine.


    NbP3d(myclass; ML: MLine) returns Integer;
    	---Purpose: Returns the number of 3d points of a MLine.


    Value(myclass; ML: MLine; U: Real; tabPt: out Array1OfPnt);
    	---Purpose: returns the 3d points of the multipoint <MPointIndex>
    	--          when only 3d points exist.


    Value(myclass; ML: MLine; U: Real; tabPt2d: out Array1OfPnt2d);
    	---Purpose: returns the 2d points of the multipoint <MPointIndex>
    	--          when only 2d points exist.


    Value(myclass; ML: MLine; U: Real; 
          tabPt: out Array1OfPnt; tabPt2d: out Array1OfPnt2d);
    	---Purpose: returns the 3d and 2d points of the multipoint 
    	--          <MPointIndex>.


    D1(myclass; ML: MLine; U: Real; tabV: out Array1OfVec)
    returns Boolean;
    	---Purpose: returns the 3d derivative values of the multipoint 
    	--          <MPointIndex> when only 3d points exist.


    D1(myclass; ML: MLine; U: Real; tabV2d: out Array1OfVec2d)
    returns Boolean;
    	---Purpose: returns the 2d derivative values of the multipoint 
    	--          <MPointIndex> only when 2d points exist.


    D1(myclass; ML: MLine; U: Real; 
             tabV: out Array1OfVec; tabV2d: out Array1OfVec2d)
    returns Boolean;
    	---Purpose: returns the 3d and 2d derivative values of the multipoint 
    	--          <MPointIndex>.


end TheLineTool;    
    
