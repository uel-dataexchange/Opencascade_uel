-- File:	RWStepShape_RWSweptFaceSolid.cdl
-- Created:	Mon Mar 15 16:13:04 1999
-- Author:	data exchange team
--		<det@androx.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class RWSweptFaceSolid from RWStepShape 

	---Purpose: Read & Write Module for SweptFaceSolid

uses

     Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SweptFaceSolid from StepShape,
     EntityIterator from Interface

is
    	Create returns RWSweptFaceSolid;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable SweptFaceSolid from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : SweptFaceSolid from StepShape);

	Share(me; ent : SweptFaceSolid from StepShape; iter : in out EntityIterator);


end RWSweptFaceSolid;
