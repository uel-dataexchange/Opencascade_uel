-- File:        BSplineCurveWithKnots.cdl
-- Created:     Fri Dec  1 11:11:14 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class BSplineCurveWithKnots from StepGeom 

inherits BSplineCurve from StepGeom 

uses

	HArray1OfInteger from TColStd, 
	HArray1OfReal from TColStd, 
	KnotType from StepGeom, 
	Integer from Standard, 
	Real from Standard, 
	HAsciiString from TCollection, 
	HArray1OfCartesianPoint from StepGeom, 
	BSplineCurveForm from StepGeom, 
	Logical from StepData
is

	Create returns mutable BSplineCurveWithKnots;
	---Purpose: Returns a BSplineCurveWithKnots


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aDegree : Integer from Standard;
	      aControlPointsList : mutable HArray1OfCartesianPoint from StepGeom;
	      aCurveForm : BSplineCurveForm from StepGeom;
	      aClosedCurve : Logical from StepData;
	      aSelfIntersect : Logical from StepData) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aDegree : Integer from Standard;
	      aControlPointsList : mutable HArray1OfCartesianPoint from StepGeom;
	      aCurveForm : BSplineCurveForm from StepGeom;
	      aClosedCurve : Logical from StepData;
	      aSelfIntersect : Logical from StepData;
	      aKnotMultiplicities : mutable HArray1OfInteger from TColStd;
	      aKnots : mutable HArray1OfReal from TColStd;
	      aKnotSpec : KnotType from StepGeom) is virtual;

	-- Specific Methods for Field Data Access --

	SetKnotMultiplicities(me : mutable; aKnotMultiplicities : mutable HArray1OfInteger);
	KnotMultiplicities (me) returns mutable HArray1OfInteger;
	KnotMultiplicitiesValue (me; num : Integer) returns Integer;
	NbKnotMultiplicities (me) returns Integer;
	SetKnots(me : mutable; aKnots : mutable HArray1OfReal);
	Knots (me) returns mutable HArray1OfReal;
	KnotsValue (me; num : Integer) returns Real;
	NbKnots (me) returns Integer;
	SetKnotSpec(me : mutable; aKnotSpec : KnotType);
	KnotSpec (me) returns KnotType;

fields

	knotMultiplicities : HArray1OfInteger from TColStd;
	knots : HArray1OfReal from TColStd;
	knotSpec : KnotType from StepGeom; -- an Enumeration

end BSplineCurveWithKnots;
