-- File:	MNaming_NamingRetrievalDriver.cdl
-- Created:	Wed Sep 17 17:08:38 1997
-- Author:	Isabelle GRIGNON
--		<isg@bigbox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997

class NamingRetrievalDriver from MNaming inherits ARDriver from MDF

	---Purpose: 

uses RRelocationTable from MDF,
     Attribute        from PDF,
     Attribute        from TDF, 
     MessageDriver    from CDM

is


    Create(theMessageDriver : MessageDriver from CDM)  -- Version 0
    returns mutable NamingRetrievalDriver from MNaming;
    

    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type: Constraint from PDataStd.

    NewEmpty (me)  returns mutable Attribute from TDF;


    Paste(me;
    	  Source     :         Attribute from PDF;
    	  Target     : mutable Attribute from TDF;
    	  RelocTable : RRelocationTable  from MDF);


end NamingRetrievalDriver;
