-- File:	PrsMgr_ModedPresentation.cdl
-- Created:	Mon Jan 30 17:56:50 1995
-- Author:	Mister rmi
--		<rmi@pernox>
---Copyright:	 Matra Datavision 1995

class ModedPresentation from PrsMgr

uses
    Presentation from PrsMgr

is
    Create 
    returns  ModedPresentation from PrsMgr;
    
    Create(aPresentation:Presentation from PrsMgr;
           aMode: Integer from Standard) 
    returns  ModedPresentation from PrsMgr;
    
    Presentation(me) returns Presentation from PrsMgr
    is static;

    Mode(me) returns Integer from Standard;

    
fields

    myPresentation: Presentation from PrsMgr;
    myMode: Integer from Standard;
    
end ModedPresentation from PrsMgr;
    
