-- File:	IGESSolid_ToolSphericalSurface.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolSphericalSurface  from IGESSolid

    ---Purpose : Tool to work on a SphericalSurface. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses SphericalSurface from IGESSolid,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolSphericalSurface;
    ---Purpose : Returns a ToolSphericalSurface, ready to work


    ReadOwnParams (me; ent : mutable SphericalSurface;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : SphericalSurface;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : SphericalSurface;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a SphericalSurface <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : SphericalSurface) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : SphericalSurface;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : SphericalSurface; entto : mutable SphericalSurface;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : SphericalSurface;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolSphericalSurface;
