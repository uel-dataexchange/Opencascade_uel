-- File:	TDF_DeltaOnForget.cdl
--      	---------------------
-- Author:	DAUTRY Philippe
--		<fid@fox.paris1.matra-dtv.fr>
---Copyright:	 MATRA DATAVISION 1997

---Version:	0.0
---History:	Version	Date		Purpose
--		0.0	Nov  3 1997	Creation
--		1.0	Jul  6 1998	Separation Forget/Resume

class DeltaOnForget from TDF inherits AttributeDelta from TDF

	---Purpose: This class provides default services for an
	--          AttributeDelta on an Forget action.
	--          
	--          Applying this AttributeDelta means RESUMING its
	--          attribute.

uses

    Attribute from TDF

is

    Create(anAtt : Attribute from TDF)
    	returns mutable DeltaOnForget from TDF;
	---Purpose: Creates a TDF_DeltaOnForget.

    Apply (me : mutable)
    	is redefined static;
    	---Purpose: Applies the delta to the attribute.

end DeltaOnForget;
