-- File:        GeometricSet.cdl
-- Created:     Fri Dec  1 11:11:21 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class GeometricSet from StepShape 

inherits GeometricRepresentationItem from StepGeom

uses

	HArray1OfGeometricSetSelect from StepShape, 
	GeometricSetSelect from StepShape, 
	HAsciiString from TCollection
is

	Create returns mutable GeometricSet;
	---Purpose: Returns a GeometricSet


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aElements : mutable HArray1OfGeometricSetSelect from StepShape) is virtual;

	-- Specific Methods for Field Data Access --

	SetElements(me : mutable; aElements : mutable HArray1OfGeometricSetSelect);
	Elements (me) returns mutable HArray1OfGeometricSetSelect;
	ElementsValue (me; num : Integer) returns GeometricSetSelect;
	NbElements (me) returns Integer;

fields

	elements : HArray1OfGeometricSetSelect from StepShape; -- a SelectType

end GeometricSet;
