-- File:	StepFEA_ElementOrElementGroup.cdl
-- Created:	Tue Feb  4 10:39:08 2003 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class ElementOrElementGroup from StepFEA
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type ElementOrElementGroup

uses
    ElementRepresentation from StepFEA,
    ElementGroup from StepFEA

is
    Create returns ElementOrElementGroup from StepFEA;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of ElementOrElementGroup select type
	--          1 -> ElementRepresentation from StepFEA
	--          2 -> ElementGroup from StepFEA
	--          0 else

    ElementRepresentation (me) returns ElementRepresentation from StepFEA;
	---Purpose: Returns Value as ElementRepresentation (or Null if another type)

    ElementGroup (me) returns ElementGroup from StepFEA;
	---Purpose: Returns Value as ElementGroup (or Null if another type)

end ElementOrElementGroup;
