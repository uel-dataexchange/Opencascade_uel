-- File:        StyleContextSelect.cdl
-- Created:     Fri Dec  1 11:11:11 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class StyleContextSelect from StepVisual inherits SelectType from StepData

	-- <StyleContextSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : Representation, RepresentationItem, PresentationSet

uses

	Representation from StepRepr,
	RepresentationItem from StepRepr,
	PresentationSet from StepVisual
is

	Create returns StyleContextSelect;
	---Purpose : Returns a StyleContextSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a StyleContextSelect Kind Entity that is :
	--        1 -> Representation
	--        2 -> RepresentationItem
	--        3 -> PresentationSet
	--        0 else

	Representation (me) returns any Representation;
	---Purpose : returns Value as a Representation (Null if another type)

	RepresentationItem (me) returns any RepresentationItem;
	---Purpose : returns Value as a RepresentationItem (Null if another type)

	PresentationSet (me) returns any PresentationSet;
	---Purpose : returns Value as a PresentationSet (Null if another type)


end StyleContextSelect;

