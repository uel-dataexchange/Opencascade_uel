-- File:      BlendFunc_CSCircular.cdl
-- Created:   Wed Jan  4 10:32:38 1995
-- Author:    Jacques GOUSSARD
---Copyright: Matra Datavision 1995


class CSCircular from BlendFunc

inherits CSFunction from Blend

	---Purpose: 

uses Vector          from math,
     Matrix          from math,
     Ax1             from gp,
     Vec             from gp,
     Vec2d           from gp,
     Pnt             from gp,
     Pnt2d           from gp,
     Circ            from gp,
     Array1OfPnt     from TColgp,
     Array1OfVec     from TColgp,
     Array1OfPnt2d   from TColgp,
     Array1OfVec2d   from TColgp,
     Array1OfReal    from TColStd,
     Array1OfInteger from TColStd,
     Shape           from GeomAbs,
     Point           from Blend,
     SectionShape    from BlendFunc,
     ParameterisationType from Convert,
     HCurve          from Adaptor3d,
     HSurface        from Adaptor3d,
     Function        from Law

is

    Create(S: HSurface from Adaptor3d; C: HCurve from Adaptor3d; CGuide: HCurve from Adaptor3d;
           L: Function from Law)

	---Purpose: Creates a function for a circular blending between
	--          a curve  <C> and a surface  <S>.  The direction of
	--          the planes are given by <CGuide>.  The position of
	--          the plane is  determined on  the  curve <C>.   <L>
	--          defines  the change of  parameter between  <C> and
	--          <CGuide>.  So, the planes are defined as described
	--          below :
	--          t is the current parameter on the guide line.
	--          Pguide = C(L(t)); Nguide = CGuide'(t)/||CGuide'(t)||
    
    	returns CSCircular from BlendFunc;
	

    NbVariables(me)
    
    	returns Integer from Standard
	is redefined;


    NbEquations(me)
    	---Purpose: returns the number of equations of the function (3).
    	returns Integer from Standard;

    Value(me: in out; X: Vector; F: out Vector)
    	---Purpose: computes the values <F> of the Functions for the 
    	--          variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    	returns Boolean from Standard;
    
    
    Derivatives(me: in out; X: Vector; D: out Matrix)
    	---Purpose: returns the values <D> of the derivatives for the 
    	--          variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    returns Boolean from Standard;
    
    
    Values(me: in out; X: Vector; F: out Vector; D: out Matrix)
    	---Purpose: returns the values <F> of the functions and the derivatives
    	--          <D> for the variable <X>.
    	--          Returns True if the computation was done successfully, 
    	--          False otherwise.

    returns Boolean from Standard;


    Set(me: in out; Param: Real from Standard)
    
    	;
	    
    Set(me: in out; First, Last: Real from Standard)
    ;
    

    GetTolerance(me; Tolerance: out Vector from math; Tol: Real from Standard)
    
    	;


    GetBounds(me; InfBound,SupBound: out Vector from math)
    
    	;

    IsSolution(me: in out; Sol: Vector from math; Tol: Real from Standard)
    
    	returns Boolean from Standard
    
    	;

    PointOnS(me)
    
    	returns Pnt from gp
	---C++: return const&
	;

    PointOnC(me)
    
    	returns Pnt from gp
	---C++: return const&
	;


    Pnt2d(me)
    
	---Purpose: Returns U,V coordinates of the point on the surface.
    
    	returns Pnt2d from gp
	---C++: return const&
	;


    ParameterOnC(me)
    
	---Purpose: Returns parameter of the point on the curve.

    	returns Real from Standard
	;


    IsTangencyPoint(me)
    
    	returns Boolean from Standard
	;

    TangentOnS(me)
    
    	returns Vec from gp
	---C++: return const&
	;

    Tangent2d(me)
    
    	returns Vec2d from gp
	---C++: return const&
	;

    TangentOnC(me)
    
    	returns Vec from gp
	---C++: return const&
	;


    Tangent(me; U,V: Real from Standard;
                TgS,NormS: out Vec from gp);
    
	---Purpose: Returns the tangent vector at the section,
	--          at the beginning and the end of the section, and
	--          returns the normal (of the surface) at
	--          these points.

-- methodes hors template (en plus du create)

    Set(me: in out; Radius : Real from Standard;
                    Choix: Integer from Standard)
    
    	is static;


    Set(me: in out; TypeSection: SectionShape from BlendFunc)
    	---Purpose: Sets  the  type  of   section generation   for the
    	--          approximations. 
    	is static;



    Section(me: in out; Param: Real from Standard;
                        U,V,W: Real from Standard;
                        Pdeb,Pfin: out Real from Standard;
                        C: out Circ from gp)
	
	is static;

    Section(me: in out; P: Point from Blend;
			Poles     : out Array1OfPnt   from TColgp;
			DPoles    : out Array1OfVec   from TColgp;
			D2Poles   : out Array1OfVec   from TColgp;
    	                Poles2d   : out Array1OfPnt2d from TColgp;
			DPoles2d  : out Array1OfVec2d from TColgp;
			D2Poles2d : out Array1OfVec2d from TColgp;
			Weigths   : out Array1OfReal  from TColStd;
			DWeigths  : out Array1OfReal  from TColStd;
                        D2Weigths : out Array1OfReal  from TColStd)

	---Purpose: Used for the first and last section 
	--          The method returns Standard_True if the derivatives
	--          are computed, otherwise it returns Standard_False.

    	returns Boolean from Standard

    	is redefined;    


    GetSection(me: in out; Param: Real from Standard;
                           U,V,W: Real from Standard;
		  	   tabP : out Array1OfPnt from TColgp;
			   tabV : out Array1OfVec from TColgp)

        returns Boolean from Standard
	
	is static;


--- Pour les approximations

    IsRational(me) returns Boolean
	---Purpose: Returns  if the section is rationnal
    is static;

    GetSectionSize(me) returns Real
    	---Purpose:  Returns the length of the maximum section
    is static;
    
    GetMinimalWeight(me; Weigths  : out Array1OfReal  from TColStd)
    	---Purpose: Compute the minimal value of weight for each poles
    	--          of all sections.
    is static;

    NbIntervals(me; S : Shape from GeomAbs) returns Integer
	---Purpose: Returns  the number  of  intervals for  continuity
	--          <S>. May be one if Continuity(me) >= <S>
    is static;
    
    Intervals(me; T : in out Array1OfReal from TColStd; 
    	          S : Shape from GeomAbs)
	---Purpose: Stores in <T> the  parameters bounding the intervals
	--          of continuity <S>.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
--    raises
--    	OutOfRange from Standard 
    is static;

    GetShape(me: in out;
                 NbPoles   : out Integer from Standard;
    	    	 NbKnots   : out Integer from Standard;
                 Degree    : out Integer from Standard;
                 NbPoles2d : out Integer from Standard)

    	is static;
	
    GetTolerance(me; 
    	    	 BoundTol, SurfTol, AngleTol : Real;
		 Tol3d : out Vector;
		 Tol1D : out Vector )
	---Purpose: Returns the tolerance to reach in approximation
	--          to respecte
	--          BoundTol error at the Boundary
	--          AngleTol tangent error at the Boundary
	--          SurfTol error inside the surface.
        is static;

    Knots(me: in out; TKnots: out Array1OfReal from TColStd)
    
	is static;


    Mults(me: in out; TMults: out Array1OfInteger from TColStd)
    
	is static;


    Section(me: in out ; P: Point from Blend;
                         Poles    : out Array1OfPnt   from TColgp;
		         DPoles   : out Array1OfVec   from TColgp;
  	                 Poles2d  : out Array1OfPnt2d from TColgp;
		         DPoles2d : out Array1OfVec2d from TColgp;
		         Weigths  : out Array1OfReal  from TColStd;
		         DWeigths : out Array1OfReal  from TColStd)

	---Purpose: Used for the first and last section 

    	returns Boolean from Standard

    	is static;


    Section(me: in out ; P: Point from Blend;
                         Poles    : out Array1OfPnt   from TColgp;
    	                 Poles2d  : out Array1OfPnt2d from TColgp;
		         Weigths  : out Array1OfReal  from TColStd)


    	is static;

    Resolution(me; 
    	       IC2d : Integer from Standard;
	       Tol  : Real from Standard;
	       TolU, TolV : out Real from Standard);

fields
    surf     : HSurface from Adaptor3d;
    curv     : HCurve from Adaptor3d;
    guide    : HCurve from Adaptor3d;
    law      : Function from Law;

    pts      : Pnt     from gp;
    ptc      : Pnt     from gp;
    pt2d     : Pnt2d   from gp;
    prmc     : Real    from Standard;
    dprmc    : Real    from Standard;
    istangent: Boolean from Standard;
    tgs      : Vec     from gp;
    tg2d     : Vec2d   from gp;
    tgc      : Vec     from gp;

    ray      : Real    from Standard;
    choix    : Integer from Standard;
    d1gui    : Vec     from gp;
    d2gui    : Vec     from gp;
    nplan    : Vec     from gp;
    normtg   : Real    from Standard;

    maxang   : Real    from Standard;
    minang   : Real    from Standard;    
    mySShape : SectionShape from BlendFunc;
    myTConv  : ParameterisationType from Convert;

end CSCircular;
