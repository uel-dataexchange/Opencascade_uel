-- File:        MeasureRepresentationItemAndQualifiedRepresentationItem.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWMeasureRepresentationItemAndQualifiedRepresentationItem from RWStepShape

	---Purpose : Read & Write Module for MeasureRepresentationItemAndQualifiedRepresentationItem

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     MeasureRepresentationItemAndQualifiedRepresentationItem from StepShape,
     EntityIterator from Interface

is

	Create returns RWMeasureRepresentationItemAndQualifiedRepresentationItem;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable MeasureRepresentationItemAndQualifiedRepresentationItem from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : MeasureRepresentationItemAndQualifiedRepresentationItem from StepShape);

	Share(me; ent : MeasureRepresentationItemAndQualifiedRepresentationItem from StepShape; iter : in out EntityIterator);

end RWMeasureRepresentationItemAndQualifiedRepresentationItem;
