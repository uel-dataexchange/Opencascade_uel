-- File:	IGESDefs_ToolUnitsData.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolUnitsData  from IGESDefs

    ---Purpose : Tool to work on a UnitsData. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses UnitsData from IGESDefs,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolUnitsData;
    ---Purpose : Returns a ToolUnitsData, ready to work


    ReadOwnParams (me; ent : mutable UnitsData;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : UnitsData;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : UnitsData;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a UnitsData <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : UnitsData) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : UnitsData;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : UnitsData; entto : mutable UnitsData;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : UnitsData;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolUnitsData;
