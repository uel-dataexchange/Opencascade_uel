-- File:	RWStepShape_RWAngularSize.cdl
-- Created:	Tue Apr 18 16:42:57 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWAngularSize from RWStepShape

    ---Purpose: Read & Write tool for AngularSize

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    AngularSize from StepShape

is
    Create returns RWAngularSize from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : AngularSize from StepShape);
	---Purpose: Reads AngularSize

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: AngularSize from StepShape);
	---Purpose: Writes AngularSize

    Share (me; ent : AngularSize from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWAngularSize;
