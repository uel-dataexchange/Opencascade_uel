-- File:	IGESGraph_ToolDefinitionLevel.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolDefinitionLevel  from IGESGraph

    ---Purpose : Tool to work on a DefinitionLevel. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses DefinitionLevel from IGESGraph,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolDefinitionLevel;
    ---Purpose : Returns a ToolDefinitionLevel, ready to work


    ReadOwnParams (me; ent : mutable DefinitionLevel;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : DefinitionLevel;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : DefinitionLevel;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a DefinitionLevel <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : DefinitionLevel) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : DefinitionLevel;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : DefinitionLevel; entto : mutable DefinitionLevel;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : DefinitionLevel;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolDefinitionLevel;
