-- File:	StepFEA_SymmetricTensor22d.cdl
-- Created:	Thu Dec 12 17:51:06 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class SymmetricTensor22d from StepFEA
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type SymmetricTensor22d

uses
    HArray1OfReal from TColStd

is
    Create returns SymmetricTensor22d from StepFEA;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of SymmetricTensor22d select type
	--          1 -> HArray1OfReal from TColStd
	--          0 else

    AnisotropicSymmetricTensor22d (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns Value as AnisotropicSymmetricTensor22d (or Null if another type)

end SymmetricTensor22d;
