-- File:        AutoDesignActualDateAndTimeAssignment.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWAutoDesignActualDateAndTimeAssignment from RWStepAP214

	---Purpose : Read & Write Module for AutoDesignActualDateAndTimeAssignment

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     AutoDesignActualDateAndTimeAssignment from StepAP214,
     EntityIterator from Interface

is

	Create returns RWAutoDesignActualDateAndTimeAssignment;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable AutoDesignActualDateAndTimeAssignment from StepAP214);

	WriteStep (me; SW : in out StepWriter; ent : AutoDesignActualDateAndTimeAssignment from StepAP214);

	Share(me; ent : AutoDesignActualDateAndTimeAssignment from StepAP214; iter : in out EntityIterator);

end RWAutoDesignActualDateAndTimeAssignment;
