-- File:	LocOpe_Spliter.cdl
-- Created:	Fri Jan 12 10:57:27 1996
-- Author:	Jacques GOUSSARD
--		<jag@bravox>
---Copyright:	 Matra Datavision 1996


class Spliter from LocOpe

	---Purpose: 

uses Shape                     from TopoDS,
     Face                      from TopoDS,
     ProjectedWires            from LocOpe,
     ListOfShape               from TopTools,
     DataMapOfShapeListOfShape from TopTools



raises NotDone      from StdFail,
       NullObject   from Standard,
       NoSuchObject from Standard

is

    Create
	---Purpose: Empty constructor.
    	returns Spliter from LocOpe;
    	---C++: inline


    Create(S: Shape from TopoDS)
	---Purpose: Creates the algorithm on the shape <S>.
	---C++: inline
    	returns Spliter from LocOpe;


    Init(me: in out; S: Shape from TopoDS)
	---Purpose: Initializes the algorithm on the shape <S>.
	---C++: inline
    	is static;


    Perform(me: in out; PW: ProjectedWires from LocOpe)
			
	raises NullObject from Standard		
    	is static;


    IsDone(me)
    
	---C++: inline
    	returns Boolean from Standard
	is static;



    ResultingShape(me)
	---Purpose: Returns the new shape
    	returns Shape from TopoDS
	---C++: return const&
	---C++: inline
	raises NotDone from StdFail
	is static;
	

    Shape(me)
	---Purpose: Returns the initial shape
    	returns Shape from TopoDS
	---C++: return const&
	---C++: inline
	is static;



    DirectLeft(me)
	---Purpose: Returns  the faces   which  are the  left of   the
	--          projected wires and which are
    	returns ListOfShape from TopTools
	---C++: return const&
	raises NotDone from StdFail
	--- The exception is raised when IsDone returns <Standard_False>.
	is static;


    Left(me)
	---Purpose: Returns the faces of the "left" part on the shape.
	--          (It  is build   from  DirectLeft,  with  the faces
	--          connected to this set, and so on...).
    	returns ListOfShape from TopTools
	---C++: return const&
	raises NotDone from StdFail
	--- The exception is raised when IsDone returns <Standard_False>.
	is static;


    DescendantShapes(me: in out; S: Shape from TopoDS)
    	---Purpose: Returns the list of descendant shapes of <S>.
    	returns ListOfShape from TopTools
	---C++: return const&
	raises NotDone from StdFail,
	       NoSuchObject from Standard
	--- The  exception  NotDone   is  raised  when  IsDone returns
	--  <Standard_False>. The exception  NoSuchObject is raised if
	--  <S> is not a subshape of the original shape.
	is static;


fields

    myShape     : Shape                     from TopoDS;
    myDone      : Boolean                   from Standard;
    myRes       : Shape                     from TopoDS;
    myMap       : DataMapOfShapeListOfShape from TopTools;
    myDLeft     : ListOfShape               from TopTools;
    myLeft      : ListOfShape               from TopTools;

end Spliter;
