-- File:	StepAP203_ClassifiedItem.cdl
-- Created:	Fri Nov 26 16:26:26 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class ClassifiedItem from StepAP203
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type ClassifiedItem

uses
    ProductDefinitionFormation from StepBasic,
    AssemblyComponentUsage from StepRepr

is
    Create returns ClassifiedItem from StepAP203;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of ClassifiedItem select type
	--          1 -> ProductDefinitionFormation from StepBasic
	--          2 -> AssemblyComponentUsage from StepRepr
	--          0 else

    ProductDefinitionFormation (me) returns ProductDefinitionFormation from StepBasic;
	---Purpose: Returns Value as ProductDefinitionFormation (or Null if another type)

    AssemblyComponentUsage (me) returns AssemblyComponentUsage from StepRepr;
	---Purpose: Returns Value as AssemblyComponentUsage (or Null if another type)

end ClassifiedItem;
