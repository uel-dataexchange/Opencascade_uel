-- File:	StepBasic_DocumentFile.cdl
-- Created:	Thu May 11 16:38:00 2000 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class DocumentFile from StepBasic
inherits Document from StepBasic

    ---Purpose: Representation of STEP entity DocumentFile

uses
    HAsciiString from TCollection,
    DocumentType from StepBasic,
    CharacterizedObject from StepBasic

is
    Create returns DocumentFile from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aDocument_Id: HAsciiString from TCollection;
                       aDocument_Name: HAsciiString from TCollection;
                       hasDocument_Description: Boolean;
                       aDocument_Description: HAsciiString from TCollection;
                       aDocument_Kind: DocumentType from StepBasic;
                       aCharacterizedObject_Name: HAsciiString from TCollection;
                       hasCharacterizedObject_Description: Boolean;
                       aCharacterizedObject_Description: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    CharacterizedObject (me) returns CharacterizedObject from StepBasic;
	---Purpose: Returns data for supertype CharacterizedObject
    SetCharacterizedObject (me: mutable; CharacterizedObject: CharacterizedObject from StepBasic);
	---Purpose: Set data for supertype CharacterizedObject

fields
    theCharacterizedObject: CharacterizedObject from StepBasic; -- supertype

end DocumentFile;
