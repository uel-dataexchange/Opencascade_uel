--
-- File:	Aspect_GraphicDriver.cdl
-- Created:	Mardi 28 janvier 1997
-- Author:	CAL
--
---Copyright:	MatraDatavision 1997
--

deferred class GraphicDriver from Aspect inherits TShared

is

	Initialize;

end GraphicDriver from Aspect;
