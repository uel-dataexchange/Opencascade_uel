-- File:        Pcurve.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPcurve from RWStepGeom

	---Purpose : Read & Write Module for Pcurve

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Pcurve from StepGeom,
     EntityIterator from Interface

is

	Create returns RWPcurve;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Pcurve from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : Pcurve from StepGeom);

	Share(me; ent : Pcurve from StepGeom; iter : in out EntityIterator);

end RWPcurve;
