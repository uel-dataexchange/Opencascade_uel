-- File:	RWStepBasic_RWConversionBasedUnitAndAreaUnit.cdl
-- Created:	Tue Oct 12 13:47:04 1999
-- Author:	data exchange team
--		<det@friendox>
---Copyright:	 Matra Datavision 1999


class RWConversionBasedUnitAndAreaUnit from RWStepBasic 

	---Purpose: Read & Write Module for RWConversionBasedUnitAndAreaUnit

uses
    
    Check from Interface,
    StepReaderData from StepData,
    StepWriter from StepData,
    ConversionBasedUnitAndAreaUnit from StepBasic,
    EntityIterator from Interface

is

    Create returns RWConversionBasedUnitAndAreaUnit from RWStepBasic;
    
    ReadStep (me; data: StepReaderData; num : Integer;
	          ach : in out Check; ent : mutable ConversionBasedUnitAndAreaUnit from StepBasic);

    WriteStep (me; SW : in out StepWriter; ent : ConversionBasedUnitAndAreaUnit from StepBasic);

    Share(me; ent : ConversionBasedUnitAndAreaUnit from StepBasic; iter : in out EntityIterator);
    
end RWConversionBasedUnitAndAreaUnit;
