-- File:	RWStepRepr_RWStructuralResponsePropertyDefinitionRepresentation.cdl
-- Created:	Sun Dec 15 10:59:25 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWStructuralResponsePropertyDefinitionRepresentation from RWStepRepr

    ---Purpose: Read & Write tool for StructuralResponsePropertyDefinitionRepresentation

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    StructuralResponsePropertyDefinitionRepresentation from StepRepr

is
    Create returns RWStructuralResponsePropertyDefinitionRepresentation from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : StructuralResponsePropertyDefinitionRepresentation from StepRepr);
	---Purpose: Reads StructuralResponsePropertyDefinitionRepresentation

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: StructuralResponsePropertyDefinitionRepresentation from StepRepr);
	---Purpose: Writes StructuralResponsePropertyDefinitionRepresentation

    Share (me; ent : StructuralResponsePropertyDefinitionRepresentation from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWStructuralResponsePropertyDefinitionRepresentation;
