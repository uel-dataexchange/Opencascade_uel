
-- File:	Graphic2d_Image.cdl
-- Created:	Tue Jun 22 16:36:51 1993
-- Author:	Jean Louis FRENKEL, Gerard GRAS
--		<jlf@stylox>
-- Modified: TCL G002A, 28-11-00, new section "inquire methods"

---Copyright:	 Matra Datavision 1993

class Image from Graphic2d inherits Primitive from Graphic2d

	---Version:

	---Purpose: This class defines the primitive Image

	---Keywords: Primitive, Image
	---Warning:
	---References:

uses
	Drawer          from Graphic2d,
	Image		from Image,
	GraphicObject	from Graphic2d,
	Length          from Quantity,
	CardinalPoints  from Aspect, 
	FStream         from Aspect,
	IFStream	from Aspect


is
	-------------------------
	-- Category: Constructors
	-------------------------

	Create (aGraphicObject: GraphicObject from Graphic2d;
		anImage: Image from Image;
		X, Y: Length from Quantity;
		adx:  Length from Quantity = 0.0;
		ady:  Length from Quantity = 0.0;
		aTypeOfPlacement: CardinalPoints
				from Aspect = Aspect_CP_Center)
	returns mutable Image from Graphic2d;
	---Level: Public
	---Purpose: Defines an image with its center location;
	--	    <X>, <Y> defines the position in the space model.
	--	    <adx>, <ady> defines an offset in the device space.
	--	    The image will be placed at this offset
	--	    according to the type of placement.
	--
	--	    CardinalPoints values :
	--		- CP_North
	--		- CP_NorthEast
	--		- CP_East
	--		- CP_SouthEast
	--		- CP_South
	--		- CP_SouthWest
	--		- CP_West
	--		- CP_NorthWest
	--		- CP_Center
	---Category: Constructors

	--------------------------
	-- Category: Draw and Pick
	--------------------------

	Draw (me : mutable; aDrawer: Drawer from Graphic2d)
	is static protected;
	---Level: Internal
	---Purpose: Draws the image at the required center location
	--	    defined by the SetCenter method.

	Pick (me : mutable;
		X, Y: ShortReal from Standard;
		aPrecision: ShortReal from Standard;
		aDrawer: Drawer from Graphic2d)
	returns Boolean from Standard is static protected;
	---Purpose: Returns Standard_True if the image <me> is picked,
	--          Standard_False if not.

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetCenter (me: mutable;
		X, Y: Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Modifies the center location of the image <me>.
	---Category: Methods to modify the class definition

	SetOffset (me: mutable;
		dx, dy: Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Modifies the offset of the image <me>.
	---Category: Methods to modify the class definition

	SetPlacement (me: mutable; aPlacement: CardinalPoints from Aspect)
	is  static;
	---Level: Public
	---Purpose: Modifies the type of placement of the image <me>.
	--
	--	    CardinalPoints values :
	--		- CP_North
	--		- CP_NorthEast
	--		- CP_East
	--		- CP_SouthEast
	--		- CP_South
	--		- CP_SouthWest
	--		- CP_West
	--		- CP_NorthWest
	--		- CP_Center
	---Category: Methods to modify the class definition

	Translate (me: mutable;
	           DX, DY: Length from Quantity) is static;
	---Level: Public
	---Purpose: Modifies the center location of the image <me>
	--          by translating it.
	---Category: Methods to modify the class definition

	Clear (me: mutable) is static;
	---Level: Public
	---Purpose: Clear the reference to this image if something
	-- 	   inside have changed,Forced the reload of this at Draw()
	--	   time.
	---Category: Methods to modify the class definition

	-------------------------------------------------------
	-- Category: Methods to manage the filling of the image
	-------------------------------------------------------

	SetSmallSize (myclass; aSize: Integer from Standard);
	---Level: Internal
	---Purpose: Defines the limit between a large image and a
	--	    small image.
	--  Warning: A small image have Height*Width <= SmallSize ().
	--	    Default 4096 = 64*64
	---Category: Methods to manage the filling of the image

	SmallSize (myclass)
	returns Integer from Standard;
	---Level: Internal
	---Purpose: Returns the limit between a large image and a
	--	    small image.
	--  Warning: A small image have Height*Width <= SmallSize ().
	---Category: Methods to manage the filling of the image

    --------------------------------------
	-- Category: Inquire methods
	--------------------------------------

    Position( me; X, Y: out Length from Quantity );  
	---Level: Public
	---Purpose: returns the position in the space model
	
	Offset( me; aX, aY: out Length from Quantity );
	---Level: Public
	---Purpose: returns the offset in the device space
	
    Placement( me ) returns CardinalPoints from Aspect;
	---Level: Public
	---Purpose: returns the type of placement
	
	Image( me ) returns Image from Image;
	---Level: Public
	---Purpose: returns the image
	
	----------------------------
	-- Category: Private methods
	----------------------------

	FillAndDraw (me; aDrawer: Drawer from Graphic2d)
	is static private;
	---Level: Internal
	---Purpose: Fills the image <me> in the drawer <aDrawer>.
	---Category: Private methods

	ComputeCenter (me;
		aDrawer: Drawer from Graphic2d;
		cx, cy: out ShortReal from  Standard)
	is static private;
	---Level: Internal
	---Purpose: Evaluates the center of the image in the device space.
	--	    Called by the methods Graphic2d_Image::Draw,
	--	    Graphic2d_Image::Pick and Graphic2d_Image::FillAndDraw.
	---Category: Private methods

	----------------------------------------------------------------------

	Save( me; aFStream: in out FStream from Aspect ) is virtual;
--	Retrieve( me; aIFStream: in out IFStream from AIS2D ) is virtual;

fields

	myImage:	  Image from Image;
	myX, myY:	  ShortReal from Standard;
	mydx, mydy:	  ShortReal from Standard;
	myPlacement:  CardinalPoints from Aspect;
	myIsModified: Boolean from Standard;

end Image from Graphic2d;
