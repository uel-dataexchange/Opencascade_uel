
-- File:	Graphic2d_Vertex.cdl
-- Created:	Mercredi 11 Aout 1993
-- Author:	CAL
--
---Copyright:	MatraDatavision 1993
--

class Vertex from Graphic2d

	---Version:

	---Purpose: This class allows the creation and update of a
	--	    2D point.

	---Keywords: Vertex, Coordinate, Point
	---Warning:
	---References:

uses
	Drawer	from Graphic2d,
	Length	from Quantity

is
	-------------------------
	-- Category: Constructors
	-------------------------

	Create
	returns Vertex from Graphic2d;
	---Level: Public
	---Purpose: Creates a point with 0.0, 0.0 coordinates.

	Create (AX, AY: Real from Standard)
	returns Vertex from Graphic2d;
	---Level: Public
	---Purpose: Creates a point with <AX>, <AY> coordinates.

	Create (AX, AY: ShortReal from Standard)
	returns Vertex from Graphic2d;
	---Level: Public
	---Purpose: Creates a point with <AX>, <AY> coordinates.

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetCoord (me: in out;
		  Xnew, Ynew: Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Modifies the coordinates of the point <me>.
	---Category: Methods to modify the class definition

	SetXCoord (me: in out;
		   Xnew: Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Modifies the X coordinate of the point <me>.
	---Category: Methods to modify the class definition

	SetYCoord (me: in out;
		   Ynew: Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Modifies the Y coordinate of the point <me>.
	---Category: Methods to modify the class definition

	----------------------------
	-- Category: Inquire methods
	----------------------------

	Coord (me;
		AX, AY: out Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Returns the coordinates of the point <me>.
	---Category: Inquire methods

	X (me) returns Length from Quantity
	is static;
	---Level: Public
	---Purpose: Returns the X coordinates of the point <me>.
	---Category: Inquire methods

	Y (me) returns Length from Quantity
	is static;
	---Level: Public
	---Purpose: Returns the Y coordinate of the point <me>.
	---Category: Inquire methods

   	IsEqual (me ; other : Vertex) returns Boolean
   	is static;
   	---Level: Public
   	---Purpose: Test if <me> and <other> are the the same vertex.
   	---C++: alias operator ==

	--------------------------
	-- Category: Class methods
	--------------------------

	Distance (myclass;
		   AV1, AV2: Vertex from Graphic2d)
	returns Length from Quantity;
	---Level: Public
	---Purpose: Returns the distance between <AV1> and <AV2>.
	---Category: Class methods

fields
	myX:	ShortReal from Standard;
	myY:	ShortReal from Standard;

end Vertex from Graphic2d;
