-- File:	IGESBasic_ToolExternalReferenceFile.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolExternalReferenceFile  from IGESBasic

    ---Purpose : Tool to work on a ExternalReferenceFile. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses ExternalReferenceFile from IGESBasic,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolExternalReferenceFile;
    ---Purpose : Returns a ToolExternalReferenceFile, ready to work


    ReadOwnParams (me; ent : mutable ExternalReferenceFile;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : ExternalReferenceFile;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : ExternalReferenceFile;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a ExternalReferenceFile <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : ExternalReferenceFile) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : ExternalReferenceFile;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : ExternalReferenceFile; entto : mutable ExternalReferenceFile;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : ExternalReferenceFile;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolExternalReferenceFile;
