-- File:	PTopoDS_Vertex.cdl
-- Created:	Wed May  5 16:53:16 1993
-- Author:	Remi LEQUETTE
--		<rle@sdsun1>
---Copyright:	 Matra Datavision 1993


class Vertex from PTopoDS inherits HShape from PTopoDS

is
    Create returns mutable Vertex from PTopoDS;
    	---Level: Internal 

end Vertex;
