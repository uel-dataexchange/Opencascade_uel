-- File:        TextStyle.cdl
-- Created:     Mon Dec  4 12:02:32 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWTextStyle from RWStepVisual

	---Purpose : Read & Write Module for TextStyle

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     TextStyle from StepVisual,
     EntityIterator from Interface

is

	Create returns RWTextStyle;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable TextStyle from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : TextStyle from StepVisual);

	Share(me; ent : TextStyle from StepVisual; iter : in out EntityIterator);

end RWTextStyle;
