-- File:	XmlMXCAFDoc_DimTolToolDriver.cdl
-- Created:	Wed Dec 10 15:02:13 2008
-- Author:	Pavel TELKOV
--		<ptv@valenox>
---Copyright:	 Open CASCADE 2008

class DimTolToolDriver from XmlMXCAFDoc  inherits ADriver from XmlMDF

        ---Purpose: Attribute Driver.

uses
    SRelocationTable from XmlObjMgt,
    RRelocationTable from XmlObjMgt,
    Persistent       from XmlObjMgt,
    MessageDriver    from CDM,
    Attribute        from TDF

is
    Create (theMsgDriver:MessageDriver from CDM)
    returns mutable DimTolToolDriver from XmlMXCAFDoc;

    NewEmpty (me)  
    returns mutable Attribute from TDF
    is redefined;

    Paste(me; theSource     : Persistent from XmlObjMgt;
              theTarget     : mutable Attribute from TDF;
              theRelocTable : out RRelocationTable from XmlObjMgt)
    returns Boolean from Standard
    is redefined;

    Paste(me; theSource     : Attribute from TDF;
              theTarget     : in out Persistent from XmlObjMgt;
              theRelocTable : out SRelocationTable from XmlObjMgt)
    is redefined;

end;
