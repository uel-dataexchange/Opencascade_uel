-- File:	VrmlConverter_DeflectionCurve.cdl
-- Created:	Tue Apr 29 14:15:41 1997
-- Author:	Alexander BRIVIN
--		<brivin@minox.nizhny.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


class DeflectionCurve from VrmlConverter 

    	---Purpose: DeflectionCurve    -  computes the presentation of
    	--          objects to be seen as  curves,   converts this  one into
    	--          VRML    objects    and    writes (adds)  into
    	--          anOStream.     All  requested properties  of   the
    	--          representation  are specify in  aDrawer.   
	--          This  kind of the presentation
    	--          is converted into IndexedLineSet ( VRML ).
        --          The computation will be made according to a maximal
        --          chordial deviation. 

uses
 
    Length       from Quantity,
    Curve        from Adaptor3d,
    Drawer       from VrmlConverter

is

    Add(myclass; anOStream: in out OStream from Standard; 
    	    	 aCurve       : in out Curve        from Adaptor3d;
    	    	 aDrawer      : Drawer       from VrmlConverter);

    ---Purpose: adds to the OStream the drawing of the curve aCurve with  
    --          respect to the maximal chordial deviation defined
    --          by the drawer aDrawer.
    --          The aspect is defined by LineAspect in aDrawer.
    --          

 
    Add(myclass; anOStream: in out OStream from Standard; 
    	    	 aCurve       : in out Curve        from Adaptor3d;
                 U1, U2       : Real         from Standard;
    	    	 aDrawer      : Drawer       from VrmlConverter);
		    
    ---Purpose: adds to the OStream the drawing of the curve aCurve with  
    --          respect to the maximal chordial deviation defined
    --          by the drawer aDrawer.
    --          The aspect is defined by LineAspect in aDrawer.
    --          The drawing will be limited between the points of parameter
    --          U1 and U2.


    Add(myclass; anOStream: in out OStream from Standard; 
    	    	 aCurve       : in out Curve        from Adaptor3d;
    	    	 aDeflection  : Real         from Standard;
    	    	 aLimit       : Real         from Standard);

    ---Purpose: adds to the OStream the drawing of the curve aCurve with  
    --          respect to the maximal chordial deviation aDeflection.
    --          The aspect is the current aspect


    Add(myclass; anOStream:  in out OStream from Standard;
    	    	 aCurve       : in out Curve        from Adaptor3d;
    	    	 aDeflection  : Real         from Standard;
    	    	 aDrawer      : Drawer       from VrmlConverter);

    ---Purpose: adds to the OStream the drawing of the curve aCurve with  
    --          respect to the maximal chordial deviation aDeflection.
    --          The aspect is the current aspect


    Add(myclass; anOStream: in out OStream from Standard; 
    	    	 aCurve       : in out Curve        from Adaptor3d;
                 U1, U2       : Real         from Standard;
    	    	 aDeflection  : Real         from Standard);
		 
    ---Purpose: adds to the OStream the drawing of the curve aCurve with  
    --          respect to the maximal chordial deviation aDeflection.
    --          The aspect is the current aspect
    --          The drawing will be limited between the points of parameter
    --          U1 and U2.


end DeflectionCurve;
