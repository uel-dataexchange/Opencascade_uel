-- File:	MultiCurve.cdl
-- Created:	Mon Dec  2 13:52:19 1991
-- Author:	Laurent PAINNOT
--		<lpa@topsn3>
---Copyright:	 Matra Datavision 1991, 1992




class MultiCurve from AppParCurves

    	---Purpose: This class describes a MultiCurve approximating a Multiline.
    	--          As a Multiline is a set of n lines, a MultiCurve is a set 
    	--          of n curves. These curves are Bezier curves.
    	--          A MultiCurve is composed of m MultiPoint. 
    	--          The approximating degree of these n curves is the same for 
    	--          each one.
    	--
    	--
    	--   Example of a MultiCurve composed of MultiPoints:
    	-- 
    	--      P1______P2_____P3______P4________........_____PNbMPoints
    	--
    	--      Q1______Q2_____Q3______Q4________........_____QNbMPoints
    	--      .                                               .
    	--      .                                               .
    	--      .                                               .
    	--      R1______R2_____R3______R4________........_____RNbMPoints
    	--
    	--     
    	--      Pi, Qi, ..., Ri are points of dimension 2 or 3.
    	--      
    	--      (Pi, Qi, ...Ri), i= 1,...NbPoles are MultiPoints.
    	--      each MultiPoint has got NbPol Poles.


uses MultiPoint              from AppParCurves,
     HArray1OfMultiPoint     from AppParCurves,
     Array1OfMultiPoint      from AppParCurves,
     Array1OfPnt             from TColgp,
     Array1OfPnt2d           from TColgp,
     Pnt                     from gp,
     Pnt2d                   from gp,
     Vec                     from gp,
     Vec2d                   from gp,
     OStream                 from Standard
     
  
raises OutOfRange        from Standard,
       DimensionError    from Standard,
       ConstructionError from Standard

is

    Create returns MultiCurve;
    	---Purpose: returns an indefinite MultiCurve.


    Create(NbPol: Integer)
    	---Purpose: creates a MultiCurve, describing Bezier curves all 
    	--          containing the same number of MultiPoint.
    	--          An exception is raised if Degree < 0.


    returns MultiCurve from AppParCurves
    raises OutOfRange from Standard;


    Create(tabMU: Array1OfMultiPoint)
    	---Purpose: creates a MultiCurve, describing Bezier curves all 
    	--          containing the same number of MultiPoint.
    	--          Each MultiPoint must have NbCurves Poles.

    returns MultiCurve from AppParCurves
    raises ConstructionError from Standard;
    
    
    Delete(me:out) is virtual;
    ---C++: alias "Standard_EXPORT virtual ~AppParCurves_MultiCurve(){Delete();}"
    
    SetNbPoles(me: in out; nbPoles: Integer)
    	---Purpose: The number of poles of the MultiCurve 
    	--          will be set to <nbPoles>.

    is static;
    
    

    SetValue(me: in out; Index: Integer; 
    	     MPoint: MultiPoint from AppParCurves)
    	---Purpose: sets the MultiPoint of range Index to the value 
    	--          <MPoint>.
    	--          An exception is raised if Index <0 or Index >NbMPoint.

    raises OutOfRange from Standard,
    	   DimensionError from Standard
    is static;
    
    

    NbCurves(me)
    	---Purpose: Returns the number of curves resulting from the
    	-- approximation of a MultiLine.

    returns Integer
    is static;
    
    
    NbPoles(me)
    	---Purpose:  Returns the number of poles on curves resulting from the approximation of a MultiLine.
    
    returns Integer
    is virtual;
    
    
    Degree(me)
    	---Purpose: returns the degree of the curves.
    
    returns Integer
    is virtual;
    

    Dimension(me; CuIndex: Integer)
    	---Purpose: returns the dimension of the CuIndex curve.
    	--          An exception is raised if CuIndex<0 or CuIndex>NbCurves.
    returns Integer
    raises OutOfRange from Standard
    is static;
    

    Curve(me; CuIndex: Integer; TabPnt: in out Array1OfPnt)
    	---Purpose: returns the Pole array of the curve of range CuIndex.
    	--          An exception is raised if the dimension of the curve 
    	--          is 2d.

    raises OutOfRange from Standard,
    	   DimensionError from Standard
    is static;


    Curve(me; CuIndex: Integer; TabPnt: in out Array1OfPnt2d)
    	---Purpose: returns the Pole array of the curve of range CuIndex.
    	--          An exception is raised if the dimension of the curve 
    	--          is 3d.

    raises OutOfRange from Standard,
    	   DimensionError from Standard
    is static;


    Value(me; Index: Integer)
    	---Purpose: returns the Index MultiPoint. 
    	--          An exception is raised if Index <0 or Index >Degree+1.
    	---C++: return const&

    returns MultiPoint from AppParCurves
    raises OutOfRange from Standard
    is static;


    Pole(me; CuIndex, Nieme: Integer)
    	---Purpose: returns the Nieme pole of the CuIndex curve.
    	--          the curve must be a 3D curve.
    	---C++: return const&

    returns Pnt from gp
    raises OutOfRange from Standard
    is static;


    Pole2d(me; CuIndex, Nieme: Integer)
    	---Purpose: returns the Nieme pole of the CuIndex curve.
    	--          the curve must be a 2D curve.
    	---C++: return const&

    returns Pnt2d from gp
    raises OutOfRange from Standard
    is static;


    Transform(me: in out; CuIndex: Integer; x, dx, y, dy, z, dz: Real)
        ---Purpose: Applies a transformation to the curve of range 
        --          <CuIndex>.
        --          newx = x + dx*oldx
        --          newy = y + dy*oldy    for all points of the curve.
        --          newz = z + dz*oldz

    raises OutOfRange from Standard
    is static;


    Transform2d(me: in out; CuIndex: Integer; x, dx, y, dy: Real)
        ---Purpose: Applies a transformation to the Curve of range 
        --          <CuIndex>.
        --          newx = x + dx*oldx
        --          newy = y + dy*oldy    for all points of the curve.

    raises OutOfRange from Standard
    is static;


    Value(me; CuIndex: Integer; U: Real; Pt: out Pnt)
    	---Purpose: returns the value of the point with a parameter U
    	--          on the Bezier curve number CuIndex.
    	--          An exception is raised if CuIndex <0 or > NbCurves.
    	--          An exception is raised if the curve dimension is 2d.

    raises OutOfRange from Standard, 
    	   DimensionError from Standard
    is virtual;
    
    
    Value(me; CuIndex: Integer; U: Real; Pt: out Pnt2d)
    	---Purpose: returns the value of the point with a parameter U
    	--          on the Bezier curve number CuIndex.
    	--          An exception is raised if CuIndex <0 or > NbCurves.
    	--          An exception is raised if the curve dimension is 3d.

    raises OutOfRange from Standard,
    	   DimensionError from Standard
    is virtual;

    
    D1(me; CuIndex: Integer; U: Real; Pt: out Pnt; V1: out Vec)
    	---Purpose: returns the value of the point with a parameter U
    	--          on the Bezier curve number CuIndex.
    	--          An exception is raised if CuIndex <0 or > NbCurves.
    	--          An exception is raised if the curve dimension is 3d.

    raises OutOfRange from Standard,
    	   DimensionError from Standard
    is virtual;


    D1(me; CuIndex: Integer; U: Real; Pt: out Pnt2d; V1: out Vec2d)
    	---Purpose: returns the value of the point with a parameter U
    	--          on the Bezier curve number CuIndex.
    	--          An exception is raised if CuIndex <0 or > NbCurves.
    	--          An exception is raised if the curve dimension is 2d.

    raises OutOfRange from Standard,
    	   DimensionError from Standard
    is virtual;

    D2(me; CuIndex: Integer; U: Real; Pt: out Pnt; V1: out Vec; V2: out Vec)
    	---Purpose: returns the value of the point with a parameter U
    	--          on the Bezier curve number CuIndex.
    	--          An exception is raised if CuIndex <0 or > NbCurves.
    	--          An exception is raised if the curve dimension is 3d.

    raises OutOfRange from Standard,
    	   DimensionError from Standard
    is virtual;


    D2(me; CuIndex: Integer; U: Real; Pt: out Pnt2d; 
           V1: out Vec2d; V2: out Vec2d)
    	---Purpose: returns the value of the point with a parameter U
    	--          on the Bezier curve number CuIndex.
    	--          An exception is raised if CuIndex <0 or > NbCurves.
    	--          An exception is raised if the curve dimension is 2d.

    raises OutOfRange from Standard,
    	   DimensionError from Standard
    is virtual;
    

    Dump(me; o: in out OStream)
    	---Purpose: Prints on the stream o information on the current 
    	--          state of the object.
    	--          Is used to redefine the operator <<.

    is virtual;
    

fields

tabPoint:  HArray1OfMultiPoint from AppParCurves is protected;


end MultiCurve;
