-- File:	TDF.cdl
--      	--------
-- Author:	DAUTRY Philippe
--		<fid@fox.paris1.matra-dtv.fr>
---Copyright:	 MATRA DATAVISION 1997

---Version:	0.0
---History:	Version	Date		Purpose
--		0.0	Feb  5 1997	Creation


package TDF 

	---Purpose: This package provides data framework for binding
	--          features and data structures.
	--          
	--          The feature structure is a tree used to bind
	--          semantic informations about each feature together.
	--          
	--          The only one concrete   attribute defined in  this
	--           package is the TagSource attribute.This attribute
	--          is used for  random creation of child labels under
	--          a given label. Tags are randomly delivered.
  
    	---Category: GUID - AttributeID
    	--           2a96b611-ec8b-11d0-bee7-080009dc3333	TDataStd_TagSource


uses

    Standard,
    MMgt,
    TColStd,
    TCollection

is


    ---Category: DF Structure Classes
    --           ==============================================================

    class Data;
	---Purpose: The root class of this structure.

    class Label;
	---Purpose: A label is a feature in the structure.

    imported HAllocator;
    imported LabelNode;
    
    pointer LabelNodePtr to LabelNode from TDF;

    deferred class Attribute;
	---Purpose: A class each application has to implement. It is
	--          used to contain the application data.

    class TagSource;
    ---Purpose: this  attribute may be used  for automatic delivery of
    --          labels under a given label.    

    class Reference;
    ---Purpose: this  attribute is  used to  store in the  framework a
    --          reference to an other label.


    ---Category: DF Copy algorithms
    --           ==============================================================
    
    class ClosureMode;
	---Purpose:  This class provides options closure management.
    
    class ClosureTool;
	---Purpose: This class gives services around the transitive
	--          enclosure of a set of information, starting from a
	--          list of label.

    class CopyTool;
	---Purpose: This class gives services around copy/paste actions.  
	 
    class CopyLabel; 
        ---Purpose: This class gives copy of  source  label  hierarchy
	  
    class ComparisonTool;
	---Purpose: This class gives services around the comparison
	--          between two sets of information.

    ---Category: DF Transaction & Delta
    --           ==============================================================

    class Transaction;
	---Purpose: This class offers services to open, commit or
	--          abort a transaction in a more secure way than
	--          using Data from TDF.

    class Delta;
    	---Purpose: A set of AttributeDelta for a given transaction
    	--          number and reference time number.

    deferred class AttributeDelta;
    	---Purpose: Delta for a given attribute. 

    class DeltaOnAddition;
	---Purpose: Attribute delta on ADDITION action.

    class DeltaOnForget;
	---Purpose: Attribute delta on FORGET action.

    class DeltaOnResume;
	---Purpose: Attribute delta on RESUME action.

    deferred class DeltaOnRemoval;
	---Purpose: Attribute delta on REMOVAL action.

    deferred class DeltaOnModification;
	---Purpose: Attribute delta on MODIFICATION action.

    class DefaultDeltaOnRemoval;
	---Purpose: Default implementation of TDF_DeltaOnRemoval.

    class DefaultDeltaOnModification;
	---Purpose: Default implementation of TDF_DeltaOnModification.


    ---Category: DF Basic Tools
    --           ==============================================================

    class ChildIterator;
	---Purpose: A tool to iterate on the children of a label.

    class ChildIDIterator;
	---Purpose: A tool to iterate on the children of a label to
	--          find attributes with an ID.

    imported AttributeIterator;
	---Purpose: DO NOT USE THIS CLASS WITHOUT AUTHORIZATION!
    

    ---Category: DF Specific Tools
    --           ==============================================================

    class DataSet;
	---Purpose: This class is used to build a set of DF
	--          informations like labels or attributes.

    class RelocationTable;
	---Purpose: Builds a attribute relocation dictionnary useful
	--          for copy or paste actions.

    class Tool;
	---Purpose: This class provides general services.

    class LabelMapHasher;
	---Purpose: A label hasher for label maps.

    class IDFilter;
	---Purpose: This class offers filtering services around an ID list.


    ---Category: DF Classes Instantiations
    --           ==============================================================

    -- Lists
    -- -----

    class IDList instantiates List from TCollection
    	(GUID from Standard);

    class AttributeList instantiates List from TCollection
    	(Attribute from TDF);

    class LabelList instantiates List from TCollection
    	(Label from TDF);

    class AttributeDeltaList  instantiates List from TCollection
    	(AttributeDelta from TDF);

    class DeltaList instantiates List from TCollection
    	(Delta from TDF);


    -- Sequences
    -- ---------

    class AttributeSequence instantiates Sequence from TCollection
    	(Attribute from TDF);

    class LabelSequence instantiates Sequence from TCollection
    	(Label from TDF);

    -- Arrays
    -- ------

    class AttributeArray1 instantiates Array1 from TCollection
    	(Attribute from TDF);

    class HAttributeArray1 instantiates HArray1 from TCollection
    	(Attribute from TDF,
    	 AttributeArray1 from TDF);



    -- Maps
    -- ----

    class IDMap instantiates Map from TCollection
    	(GUID from Standard,
    	 GUID from Standard);

    class AttributeMap instantiates Map from TCollection
    	(Attribute from TDF,
    	 MapTransientHasher from TColStd);

    class AttributeDataMap instantiates DataMap from TCollection
    	(Attribute from TDF,
    	 Attribute from TDF,
    	 MapTransientHasher from TColStd);

    class AttributeDoubleMap instantiates DoubleMap from TCollection
    	(Attribute from TDF,
    	 Attribute from TDF,
    	 MapTransientHasher from TColStd,
    	 MapTransientHasher from TColStd);

    class AttributeIndexedMap instantiates IndexedMap from TCollection
    	(Attribute from TDF,
    	 MapTransientHasher from TColStd);


    class LabelMap instantiates Map from TCollection
    	(Label from TDF,
    	 LabelMapHasher from TDF);

    class LabelDataMap instantiates DataMap from TCollection
    	(Label from TDF,
    	 Label from TDF,
    	 LabelMapHasher from TDF);

    class LabelDoubleMap instantiates DoubleMap from TCollection
    	(Label from TDF,
    	 Label from TDF,
    	 LabelMapHasher from TDF,
    	 LabelMapHasher from TDF);

    class LabelIndexedMap instantiates IndexedMap from TCollection
    	(Label from TDF,
    	 LabelMapHasher from TDF);

    class LabelIntegerMap instantiates DataMap from TCollection
    	(Label from TDF,
	 Integer from Standard,
    	 LabelMapHasher from TDF);

    class LabelLabelMap instantiates DataMap from TCollection
    	(Label from TDF,
	 Label from TDF,
    	 LabelMapHasher from TDF);

    class GUIDProgIDMap instantiates DoubleMap from TCollection
    	(GUID from Standard,
    	 ExtendedString from TCollection,
	 GUID from Standard,
         ExtendedString from TCollection);

    ---Category: Package methods
    --           ==============================================================

    LowestID returns GUID from Standard;
	---Purpose: Returns ID "00000000-0000-0000-0000-000000000000",
	--          sometimes used as null ID.
	--          
	---C++: return const &

    UppestID returns GUID from Standard;
	---Purpose: Returns ID "ffffffff-ffff-ffff-ffff-ffffffffffff".
	--          
	---C++: return const &


    AddLinkGUIDToProgID( ID : GUID from Standard; ProgID : ExtendedString from TCollection );
      ---Purpose: Sets link between GUID and ProgID in hidden DataMap
      
    GUIDFromProgID( ProgID : ExtendedString from TCollection; ID : in out GUID from Standard )
    returns Boolean from Standard;
	---Purpose: Returns True if there is GUID for given <ProgID> then GUID is returned in <ID>
	
    
    ProgIDFromGUID( ID : GUID from Standard; ProgID : in out ExtendedString from TCollection ) 	
    returns Boolean from Standard;
	---Purpose: Returns True if there is ProgID for given <ID> then ProgID is returned in <ProgID>
    
   
end TDF;
