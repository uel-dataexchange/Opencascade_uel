-- File:	IFSelect_ModifReorder.cdl
-- Created:	Fri Mar 15 09:37:46 1996
-- Author:	Christian CAILLET
--		<cky@fidox>
---Copyright:	 Matra Datavision 1996


class ModifReorder  from IFSelect  inherits Modifier

    ---Purpose : This modifier reorders a whole model from its roots, i.e.
    --           according to <rootlast> status, it considers each of its
    --           roots, then it orders all its shared entities at any level,
    --           the result begins by the lower level entities ... ends by
    --           the roots.

uses CString, AsciiString from TCollection,
     InterfaceModel, CopyTool, Protocol from Interface, ContextModif

is

    Create (rootlast : Boolean = Standard_True) returns mutable ModifReorder;
    ---Purpose : Creates a ModifReorder. It may change the graph (it does !)
    --           If <rootlast> is True (D), roots are set at the end of packets
    --           Else, they are set at beginning (as done by AddWithRefs)

    Perform (me; ctx  : in out ContextModif;
    	     target   : mutable InterfaceModel;
    	     protocol : Protocol from Interface;
    	     TC       : in out CopyTool);
    ---Purpose : Acts by computing orders (by method All from ShareTool) then
    --           forcing them in the model. Remark that selection is ignored :
    --           ALL the model is processed in once

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns Label as "Reorder, Roots (last or first)"

fields

    thertl : Boolean;

end ModifReorder;
