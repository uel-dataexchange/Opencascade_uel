-- File:	StepAP203_CcDesignContract.cdl
-- Created:	Fri Nov 26 16:26:31 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class CcDesignContract from StepAP203
inherits ContractAssignment from StepBasic

    ---Purpose: Representation of STEP entity CcDesignContract

uses
    Contract from StepBasic,
    HArray1OfContractedItem from StepAP203

is
    Create returns CcDesignContract from StepAP203;
	---Purpose: Empty constructor

    Init (me: mutable; aContractAssignment_AssignedContract: Contract from StepBasic;
                       aItems: HArray1OfContractedItem from StepAP203);
	---Purpose: Initialize all fields (own and inherited)

    Items (me) returns HArray1OfContractedItem from StepAP203;
	---Purpose: Returns field Items
    SetItems (me: mutable; Items: HArray1OfContractedItem from StepAP203);
	---Purpose: Set field Items

fields
    theItems: HArray1OfContractedItem from StepAP203;

end CcDesignContract;
