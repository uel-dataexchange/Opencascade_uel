-- File:	TopOpeBRepDS_CurvePointInterference.cdl
-- Created:	Wed Jun 23 12:10:58 1993
-- Author:	Jean Yves LEBEY
--		<jyl@zerox>
---Copyright:	 Matra Datavision 1993


class CurvePointInterference from TopOpeBRepDS 
    inherits Interference from TopOpeBRepDS

    ---Purpose: An interference with a parameter.

uses

    Transition  from TopOpeBRepDS,
    Kind        from TopOpeBRepDS,
    OStream     from Standard    
    
is

    Create(T  : Transition from TopOpeBRepDS;
	   ST : Kind from TopOpeBRepDS;
	   S  : Integer from Standard;
	   GT : Kind from TopOpeBRepDS;
	   G  : Integer from Standard;
	   P  : Real from Standard) 
    returns mutable CurvePointInterference from TopOpeBRepDS; 
	    
    Parameter(me) returns Real from Standard
    is static;
    
    Parameter(me : mutable; P : Real from Standard)
    is static;

    Dump(me; OS : in out OStream from Standard) returns OStream
    is redefined;
    ---C++: return &
    
fields

    myParam : Real from Standard;

end CurvePointInterference from TopOpeBRepDS;
