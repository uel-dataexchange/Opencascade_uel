-- File:	StepBasic_IdentificationAssignment.cdl
-- Created:	Wed May 10 15:09:08 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class IdentificationAssignment from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity IdentificationAssignment

uses
    HAsciiString from TCollection,
    IdentificationRole from StepBasic

is
    Create returns IdentificationAssignment from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aAssignedId: HAsciiString from TCollection;
                       aRole: IdentificationRole from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    AssignedId (me) returns HAsciiString from TCollection;
	---Purpose: Returns field AssignedId
    SetAssignedId (me: mutable; AssignedId: HAsciiString from TCollection);
	---Purpose: Set field AssignedId

    Role (me) returns IdentificationRole from StepBasic;
	---Purpose: Returns field Role
    SetRole (me: mutable; Role: IdentificationRole from StepBasic);
	---Purpose: Set field Role

fields
    theAssignedId: HAsciiString from TCollection;
    theRole: IdentificationRole from StepBasic;

end IdentificationAssignment;
