-- File:	RWStepFEA_RWFeaMassDensity.cdl
-- Created:	Thu Dec 12 17:51:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFeaMassDensity from RWStepFEA

    ---Purpose: Read & Write tool for FeaMassDensity

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FeaMassDensity from StepFEA

is
    Create returns RWFeaMassDensity from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FeaMassDensity from StepFEA);
	---Purpose: Reads FeaMassDensity

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FeaMassDensity from StepFEA);
	---Purpose: Writes FeaMassDensity

    Share (me; ent : FeaMassDensity from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFeaMassDensity;
