-- File:        GlobalUncertaintyAssignedContext.cdl
-- Created:     Mon Dec  4 12:02:27 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWGlobalUncertaintyAssignedContext from RWStepRepr

	---Purpose : Read & Write Module for GlobalUncertaintyAssignedContext

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     GlobalUncertaintyAssignedContext from StepRepr,
     EntityIterator from Interface

is

	Create returns RWGlobalUncertaintyAssignedContext;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable GlobalUncertaintyAssignedContext from StepRepr);

	WriteStep (me; SW : in out StepWriter; ent : GlobalUncertaintyAssignedContext from StepRepr);

	Share(me; ent : GlobalUncertaintyAssignedContext from StepRepr; iter : in out EntityIterator);

end RWGlobalUncertaintyAssignedContext;
