-- File:	IGESDraw_ToolPerspectiveView.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolPerspectiveView  from IGESDraw

    ---Purpose : Tool to work on a PerspectiveView. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses PerspectiveView from IGESDraw,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolPerspectiveView;
    ---Purpose : Returns a ToolPerspectiveView, ready to work


    ReadOwnParams (me; ent : mutable PerspectiveView;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : PerspectiveView;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : PerspectiveView;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a PerspectiveView <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : PerspectiveView) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : PerspectiveView;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : PerspectiveView; entto : mutable PerspectiveView;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : PerspectiveView;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolPerspectiveView;
