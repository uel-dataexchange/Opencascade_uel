-- File:	Graphic3d_ArrayOfTriangles.cdl
-- Created:	04/01/01 : GG : G005 : Draw ARRAY primitives
--

class ArrayOfTriangles from Graphic3d inherits ArrayOfPrimitives from Graphic3d 

is

	-- constructor
	Create (
                maxVertexs: Integer from Standard;
		maxEdges: Integer from Standard = 0;
                hasVNormals: Boolean from Standard = Standard_False;
                hasVColors: Boolean from Standard = Standard_False;
                hasTexels: Boolean from Standard = Standard_False;
                hasEdgeInfos: Boolean from Standard = Standard_False)
	returns mutable ArrayOfTriangles from Graphic3d;
        ---Purpose: Creates an array of triangles,
        -- a triangle can be filled as:
        -- 1) creating a set of triangles defined with his vertexs.
        --    i.e:
        --    myArray = Graphic3d_ArrayOfTriangles(6)
        --    myArray->AddVertex(x1,y1,z1)
        --      ....
        --    myArray->AddVertex(x6,y6,z6)
        -- 3) creating a set of indexed triangles defined with his vertex
        --    ans edges.
        --    i.e:
        --    myArray = Graphic3d_ArrayOfTriangles(4,6)
        --    myArray->AddVertex(x1,y1,z1)
        --      ....
        --    myArray->AddVertex(x4,y4,z4)
        --    myArray->AddEdge(1)
        --    myArray->AddEdge(2)
        --    myArray->AddEdge(3)
        --    myArray->AddEdge(2)
        --    myArray->AddEdge(3)
        --    myArray->AddEdge(4)
        --
        -- <maxVertexs> defined the maximun allowed vertex number in the array.
        -- <maxEdges> defined the maximun allowed edge number in the array.
        --  Warning:
        -- When <hasVNormals> is TRUE , you must use one of
        --      AddVertex(Point,Normal)
        --  or  AddVertex(Point,Normal,Color)
        --  or  AddVertex(Point,Normal,Texel) methods.
        -- When <hasVColors> is TRUE , you must use one of
        --      AddVertex(Point,Color)
        --  or  AddVertex(Point,Normal,Color) methods.
        -- When <hasTexels> is TRUE , you must use one of
        --      AddVertex(Point,Texel)
        --  or  AddVertex(Point,Normal,Texel) methods.
        -- When <hasEdgeInfos> is TRUE , <maxEdges> must be > 0 and
        --      you must use the
        --      AddEdge(number,visibillity) method.
        --  Warning:
        -- the user is responsible about the orientation of the triangle
        -- depending of the order of the created vertex or edges and this
        -- orientation must be coherent with the vertex normal optionnaly
        -- given at each vertex (See the Orientate() methods).

end;
