-- File:        BooleanOperand.cdl
-- Created:     Fri Dec  1 11:11:10 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class BooleanOperand from StepShape 

    -- inherits SelectType from StepData

	-- <BooleanOperand> is an EXPRESS Select Type construct translation.
	-- it gathers : SolidModel, HalfSpaceSolid, CsgPrimitive, BooleanResult

uses

	SolidModel,
	HalfSpaceSolid,
	CsgPrimitive,
	BooleanResult
is

    Create returns BooleanOperand;
    ---Purpose : Returns a BooleanOperand SelectType

    SetTypeOfContent(me : in out; aTypeOfContent : Integer);

    TypeOfContent(me) returns Integer;
    	-- 1 : SolidModel,
    	-- 2 : HalfSpaceSolid,
    	-- 3 : CsgPrimitive,
    	-- 4 : BooleanResult

    SolidModel (me) returns any SolidModel;
    ---Purpose : returns Value as a SolidModel (Null if another 
    --         type)

    SetSolidModel(me : in out;
    	    	  aSolidModel : SolidModel from StepShape);

    HalfSpaceSolid (me) returns any HalfSpaceSolid;
    ---Purpose : returns Value as a HalfSpaceSolid (Null if 
    --         another type)

    SetHalfSpaceSolid(me : in out; 
    	    	      aHalfSpaceSolid : HalfSpaceSolid from StepShape);

    CsgPrimitive (me) returns CsgPrimitive;
    ---Purpose : returns Value as a CsgPrimitive (Null if another 
    --           type)
    --           CsgPrimitive is another Select Type

    SetCsgPrimitive(me : in out; 
    	    	    aCsgPrimitive : CsgPrimitive from StepShape);

    BooleanResult (me) returns any BooleanResult;
    ---Purpose : returns Value as a BooleanResult (Null if another 
    --           type)

    SetBooleanResult(me:in out;
    	    	     aBooleanResult : BooleanResult from StepShape);
    
fields

    theSolidModel     : SolidModel     from StepShape;
    theHalfSpaceSolid : HalfSpaceSolid from StepShape;
    theCsgPrimitive   : CsgPrimitive   from StepShape;  -- Select Type
    theBooleanResult  : BooleanResult  from StepShape;
    theTypeOfContent  : Integer        from Standard;

end BooleanOperand;

