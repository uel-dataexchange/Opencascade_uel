-- File:	MFunction_FunctionStorageDriver.cdl
-- Created:	Thu Jun 17 11:52:14 1999
-- Author:	Vladislav ROMASHKO
--		<vro@flox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999

class FunctionStorageDriver from MFunction inherits ASDriver from MDF

uses 
 
     SRelocationTable from MDF,
     Attribute        from TDF,
     Attribute        from PDF, 
     MessageDriver    from CDM

is 

    Create(theMessageDriver : MessageDriver from CDM)  
    returns mutable FunctionStorageDriver from MFunction;

    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;

    NewEmpty (me) returns mutable Attribute from PDF;

    Paste(me;
    	  Source     :         Attribute from TDF;
    	  Target     : mutable Attribute from PDF;
    	  RelocTable : SRelocationTable from MDF);

end FunctionStorageDriver;
