-- File:	BRepBuilderAPI_GTransform.cdl
-- Created:	Mon Dec 30 17:10:14 1996
-- Author:	Stagiaire Mary FABIEN
--		<fbi@zozox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996

class GTransform from BRepBuilderAPI inherits ModifyShape from BRepBuilderAPI

	---Purpose: Geometric transformation on a shape.
    	-- The transformation to be applied is defined as a gp_GTrsf
    	-- transformation. It may be:
    	-- -      a transformation equivalent to a gp_Trsf transformation, the
    	--    most common case: you should , however, use a BRepAPI_Transform
    	--    object to perform this kind of transformation; or
    	-- -      an affinity, or
    	-- -      more generally, any type of point transformation which may
    	--  be defined by a three row, four column matrix of transformation.
    	-- In the last two cases, the underlying geometry of the
    	-- following shapes may change:
    	-- -      a curve which supports an edge of the shape, or
    	-- -      a surface which supports a face of the shape;
    	-- For example, a circle may be transformed into an ellipse when
    	-- applying an affinity transformation.
    	-- The transformation is applied to:
    	-- -      all the curves which support edges of the shape, and
    	-- -      all the surfaces which support faces of the shape.
    	-- A GTransform object provides a framework for:
    	-- -      defining the geometric transformation to be applied,
    	-- -      implementing the transformation algorithm, and
        -- -      consulting the result.
  


uses 
    Trsf              from gp,
    GTrsf             from gp,
    Shape             from TopoDS,
    Face              from TopoDS,
    Collect           from BRepBuilderAPI,
    ShapeModification from BRepBuilderAPI,
    ListOfShape       from TopTools

-- Modified by Sergey KHROMOV - Thu Mar 27 17:45:42 2003 Begin
raises 
 NoSuchObject from Standard 
 
-- Modified by Sergey KHROMOV - Thu Mar 27 17:45:42 2003 End
is

    Create(T: GTrsf from gp)
        
    	returns GTransform from BRepBuilderAPI;
	---Purpose: Constructs a framework for applying the geometric
    	-- transformation T to a shape. Use the function
    	-- Perform to define the shape to transform.


    Create(S: Shape from TopoDS; T: GTrsf from gp; 
           Copy: Boolean from Standard  =  Standard_False)

    	returns GTransform from BRepBuilderAPI;
	---Purpose: Constructs a framework for applying the geometric
    	-- transformation T to a shape, and applies it to the shape S.
    	-- -   If the transformation T is direct and isometric (i.e. if
    	--   the determinant of the vectorial part of T is equal to
    	--   1.), and if Copy equals false (default value), the
    	--   resulting shape is the same as the original but with
    	--   a new location assigned to it.
    	-- -   In all other cases, the transformation is applied to
    	--   a duplicate of S.
    	-- Use the function Shape to access the result.
    	-- Note: the constructed framework can be reused to
    	-- apply the same geometric transformation to other
    	-- shapes: just specify them with the function Perform.


    Perform(me: in out; S   : Shape   from TopoDS; 
                        Copy: Boolean from Standard  =  Standard_False)

	---Purpose: Applies the geometric transformation defined at the
    	-- time of construction of this framework to the shape S.
    	-- -   If the transformation T is direct and isometric (i.e. if
    	--   the determinant of the vectorial part of T is equal to
    	--   1.), and if Copy equals false (default value), the
    	--   resulting shape is the same as the original but with
    	--   a new location assigned to it.
    	-- -   In all other cases, the transformation is applied to a duplicate of S.
    	--   Use the function Shape to access the result.
    	-- Note: this framework can be reused to apply the same
    	-- geometric transformation to other shapes: just specify
    	-- them by calling the function Perform again.

    	is static;

    Modified (me: in out; S : Shape from TopoDS)
    	---Purpose: Returns the list  of shapes modified from the shape
    	--          <S>. 
        ---C++: return const & 
        ---Level: Public
    returns ListOfShape from TopTools
    is redefined virtual;

-- Modified by Sergey KHROMOV - Thu Mar 27 17:43:59 2003 Begin
    ModifiedShape(me; S: Shape from TopoDS)
    	returns Shape from TopoDS
	---Purpose: Returns the modified shape corresponding to <S>.
	---C++: return const&
	raises NoSuchObject from Standard
               -- if S is not the initial shape or a sub-shape
               -- of the initial shape.
    is redefined virtual;
-- Modified by Sergey KHROMOV - Thu Mar 27 17:44:02 2003 End

fields

    myGTrsf    : GTrsf    from gp;
    myUseModif : Boolean from Standard;
    myHist     : Collect from BRepBuilderAPI;
    
end Transform;
