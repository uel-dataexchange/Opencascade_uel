-- File:	StepAP203_CertifiedItem.cdl
-- Created:	Fri Nov 26 16:26:26 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class CertifiedItem from StepAP203
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type CertifiedItem

uses
    SuppliedPartRelationship from StepRepr

is
    Create returns CertifiedItem from StepAP203;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of CertifiedItem select type
	--          1 -> SuppliedPartRelationship from StepRepr
	--          0 else

    SuppliedPartRelationship (me) returns SuppliedPartRelationship from StepRepr;
	---Purpose: Returns Value as SuppliedPartRelationship (or Null if another type)

end CertifiedItem;
