-- File:	RWStepFEA_RWGeometricNode.cdl
-- Created:	Thu Dec 12 17:51:06 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWGeometricNode from RWStepFEA

    ---Purpose: Read & Write tool for GeometricNode

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    GeometricNode from StepFEA

is
    Create returns RWGeometricNode from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : GeometricNode from StepFEA);
	---Purpose: Reads GeometricNode

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: GeometricNode from StepFEA);
	---Purpose: Writes GeometricNode

    Share (me; ent : GeometricNode from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWGeometricNode;
