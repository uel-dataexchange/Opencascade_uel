-- File:        BackgroundColour.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWBackgroundColour from RWStepVisual

	---Purpose : Read & Write Module for BackgroundColour

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     BackgroundColour from StepVisual,
     EntityIterator from Interface

is

	Create returns RWBackgroundColour;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable BackgroundColour from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : BackgroundColour from StepVisual);

	Share(me; ent : BackgroundColour from StepVisual; iter : in out EntityIterator);

end RWBackgroundColour;
