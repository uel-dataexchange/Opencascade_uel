-- File:	XSControl_Reader.cdl
-- Created:	Wed May 14 14:32:43 1997
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


class Reader  from XSControl

    	---Purpose : 
    	-- A groundwork to convert a shape to data which complies
    	-- with a particular norm. This data can be that of a whole
    	-- model or that of a specific list of entities in the model.
    	-- You specify the list using a single selection or a
    	-- combination of selections. A selection is an operator which
    	-- computes a list of entities from a list given in input. To
    	-- specify the input, you can use:
    	-- - A predefined selection such as "xst-transferrable-roots"
    	-- - A filter based on a  signature.
    	-- A signature is an operator which returns a string from an
    	-- entity according to its type.
    	-- For example:
    	-- - "xst-type" (CDL)
    	-- - "iges-level"
    	-- - "step-type".
    	-- A filter can be based on a signature by giving a value to
    	-- be matched by the string returned. For example,
    	-- "xst-type(Curve)".
    	-- If no list is specified, the selection computes its list of
    	-- entities from the whole model. To use this class, you have to
    	-- initialize the transfer norm first, as shown in the example below.
    	-- Example:
    	-- Control_Reader reader;
    	-- IFSelect_ReturnStatus status = reader.ReadFile (filename.);
    	-- When using IGESControl_Reader or STEPControl_Reader - as the
    	-- above example shows - the reader initializes the norm directly.
    	-- Note that loading the file only stores the data. It does
    	-- not translate this data. Shapes are accumulated by
    	-- successive transfers. The last shape is cleared by:
    	-- - ClearShapes which allows you to handle a new batch
    	-- - TransferRoots which restarts the list of shapes from scratch.

uses CString, OStream, Transient,
     SequenceOfTransient from TColStd, HSequenceOfTransient from TColStd,
     InterfaceModel from Interface, WorkSession from XSControl,
     ReturnStatus from IFSelect, PrintCount from IFSelect,
     Shape from TopoDS, SequenceOfShape from TopTools

is

    Create returns Reader;
    ---Purpose : Creates a Reader from scratch (creates an empty WorkSession)
    --           A WorkSession or a Controller must be provided before running

    Create (norm : CString) returns Reader;
    ---Purpose : Creates a Reader from scratch, with a norm name which
    --           identifies a Controller

    Create (WS : mutable WorkSession from XSControl;
    	    	 scratch : Boolean = Standard_True) returns Reader;
    ---Purpose : Creates a Reader from an already existing Session, with a
    --           Controller already set

    ---Purpose: Virtual destructor 
    ---C++ : alias "Standard_EXPORT virtual ~XSControl_Reader() {}"

    SetNorm (me : in out; norm : CString) returns Boolean;
    ---Purpose : Sets a specific norm to <me>
    --           Returns True if done, False if <norm> is not available

    SetWS (me : in out; WS : mutable WorkSession from XSControl;
    	    	 scratch : Boolean = Standard_True);
    ---Purpose : Sets a specific session to <me>

    WS (me) returns WorkSession from XSControl;
    ---Purpose : Returns the session used in <me>


    ReadFile (me : in out; filename : CString) returns ReturnStatus;
    ---Purpose : Loads a file and returns the read status
    --           Zero for a Model which compies with the Controller

    Model (me) returns InterfaceModel;
    ---Purpose : Returns the model. It can then be consulted (header, product)

    GiveList (me : in out; first, second : CString = "")
    	returns HSequenceOfTransient from TColStd;
    	---Purpose : Returns a list of entities from the IGES or STEP file 
    	-- according to the following rules:
    	-- - if first and second are empty strings, the whole file is selected.
    	-- - if first is an entity number or label, the entity referred to is selected.
    	-- - if first is a list of entity numbers/labels separated by commas, the entities referred to are selected,
    	-- - if first is the name of a selection in the worksession and second is not defined,
    	-- the list contains the standard output for that selection.
    	-- - if first is the name of a selection and second is defined, the criterion defined
    	-- by second is applied to the result of the first selection.
    	--  A selection is an operator which computes a list of entities from a list given in
    	-- input according to its type. If no list is specified, the selection computes its
    	-- list of entities from the whole model.
    	--   A selection can be:
    	-- - A predefined selection (xst-transferrable-mode)
    	-- - A filter based on a signature
    	-- A Signature is an operator which returns a string from an entity according to its type. For example:
    	-- - "xst-type" (CDL)
    	-- - "iges-level"
    	-- - "step-type".
    	-- For example, if you wanted to select only the advanced_faces in a STEP file you
    	-- would use the following code:
    	-- Example
    	-- Reader.GiveList("xst-transferrable-roots","step-type(ADVANCED_FACE)");
    	-- Warning
    	-- If the value given to second is incorrect, it will simply be ignored.

    GiveList (me : in out; first : CString; ent : Transient)
    	returns HSequenceOfTransient from TColStd;
    ---Purpose : Computes a List of entities from the model as follows
    --           <first> beeing a Selection, <ent> beeing an entity or a list
    --           of entities (as a HSequenceOfTransient) :
    --             the standard result of this selection applied to this list
    --           if <first> is erroneous, a null handle is returned


    NbRootsForTransfer (me : in out) returns Integer is virtual ;
    ---Purpose : Determines the list of root entities which are candidate for
    --           a transfer to a Shape, and returns the number
    --           of entities in the list

    RootForTransfer (me : in out; num : Integer = 1) returns Transient;
    ---Purpose : Returns an IGES or STEP root
    --           entity for translation. The entity is identified by its
    --           rank in a list.

    TransferOneRoot (me : in out; num : Integer = 1) returns Boolean ;
    ---Purpose : Translates a root identified by the rank num in the model.
    --           false is returned if no shape is produced.
    
    TransferOne  (me : in out; num : Integer) returns Boolean;
    ---Purpose : Translates an IGES or STEP
    --           entity identified by the rank num in the model.
    --           false is returned if no shape is produced.

    TransferEntity (me : in out; start : Transient) returns Boolean;
    ---Purpose : Translates an IGES or STEP
    --           entity in the model. true is returned if a shape is
    --           produced; otherwise, false is returned.

    TransferList (me : in out; list : HSequenceOfTransient from TColStd)
    	returns Integer;
    ---Purpose : Translates a list of entities.
    --           Returns the number of IGES or STEP entities that were
    --           successfully translated. The list can be produced with GiveList.
    --           Warning - This function does not clear the existing output shapes.

    TransferRoots (me : in out) returns Integer;
    ---Purpose : Translates all translatable
    --           roots and returns the number of successful translations.
    --           Warning - This function clears existing output shapes first.


    ClearShapes (me : in out);
    ---Purpose : Clears the list of shapes that
    --           may have accumulated in calls to TransferOne or TransferRoot.C

    NbShapes (me) returns Integer;
    ---Purpose : Returns the number of shapes produced by translation.

    Shapes (me: in out) returns SequenceOfShape from TopTools is protected;
    ---Purpose : Returns a sequence of produced shapes
    ---C++: return &
    
    Shape (me; num : Integer = 1) returns Shape from TopoDS;
    	---Purpose : Returns the shape resulting
    	-- from a translation and identified by the rank num.
    	-- num equals 1 by default. In other words, the first shape
    	-- resulting from the translation is returned.

    OneShape (me) returns Shape from TopoDS;
    	---Purpose : Returns all of the results in
    	-- a single shape which is:
    	-- - a null shape if there are no results,
    	-- - a shape if there is one result,
    	-- - a compound containing the resulting shapes if there are more than one.

    PrintCheckLoad (me; failsonly : Boolean; mode : PrintCount);
    ---Purpose : Prints the check list attached to loaded data, on the Standard
    --            Trace File (starts at cout)
    --           All messages or fails only, according to <failsonly>
    --           mode = 0 : per entity, prints messages
    --           mode = 1 : per message, just gives count of entities per check
    --           mode = 2 : also gives entity numbers

    PrintCheckTransfer (me; failsonly : Boolean; mode : PrintCount);
    	---Purpose : Displays check results for the
    	-- last translation of IGES or STEP entities to Open CASCADE
    	-- entities. Only fail messages are displayed if failsonly is
    	-- true. All messages are displayed if failsonly is
    	-- false. mode determines the contents and the order of the
    	-- messages according to the terms of the IFSelect_PrintCount enumeration.

    PrintStatsTransfer (me; what : Integer; mode : Integer = 0);
    	---Purpose :  Displays the statistics for
    	-- the last translation. what defines the kind of
    	-- statistics that are displayed as follows:
    	-- - 0 gives general statistics (number of translated roots,
    	-- number of warnings, number of fail messages),
    	-- - 1 gives root results,
    	--    - 2 gives statistics for all checked entities,
    	-- - 3 gives the list of translated entities,
    	-- - 4 gives warning and fail messages,
    	-- - 5 gives fail messages only.
    	-- The use of mode depends on the value of what. If what is 0,
    	-- mode is ignored. If what is 1, 2 or 3, mode defines the following:
    	-- - 0 lists the numbers of IGES or STEP entities in the respective model
    	-- - 1 gives the number, identifier, type and result
    	-- type for each IGES or STEP entity and/or its status
    	-- (fail, warning, etc.)
    	-- - 2 gives maximum information for each IGES or STEP entity (i.e. checks)
    	-- - 3 gives the number of entities per type of IGES or STEP entity
    	-- - 4 gives the number of IGES or STEP entities per result type and/or status
    	-- - 5 gives the number of pairs (IGES or STEP or result type and status)
    	-- - 6 gives the number of pairs (IGES or STEP or result type
    	-- and status) AND the list of entity numbers in the IGES or STEP model.
    	--   If what is 4 or 5, mode defines the warning and fail
    	-- messages as follows:
    	-- - if mode is 0 all warnings and checks per entity are returned
    	-- - if mode is 2 the list of entities per warning is returned.
    	--   If mode is not set, only the list of all entities per warning is given.
    
    GetStatsTransfer (me; list: HSequenceOfTransient from TColStd;
    	    	    	  nbMapped    : out Integer;
			  nbWithResult: out Integer;
			  nbWithFail  : out Integer);
    	---Purpose: Gives statistics about Transfer

fields

    thesession : WorkSession from XSControl;
    therootsta : Boolean is protected;              -- are roots determined
    theroots   : SequenceOfTransient is protected;  -- only roots available for Transfer
    theshapes  : SequenceOfShape;

end Reader;
