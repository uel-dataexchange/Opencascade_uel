-- File:        AutoDesignApprovalAssignment.cdl
-- Created:     Fri Dec  1 11:11:13 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class AutoDesignApprovalAssignment from StepAP214 

inherits ApprovalAssignment from StepBasic 

uses

	HArray1OfAutoDesignGeneralOrgItem from StepAP214, 
	AutoDesignGeneralOrgItem from StepAP214, 
	Approval from StepBasic
is

	Create returns mutable AutoDesignApprovalAssignment;
	---Purpose: Returns a AutoDesignApprovalAssignment


	Init (me : mutable;
	      aAssignedApproval : mutable Approval from StepBasic) is redefined;

	Init (me : mutable;
	      aAssignedApproval : mutable Approval from StepBasic;
	      aItems : mutable HArray1OfAutoDesignGeneralOrgItem from StepAP214) is virtual;

	-- Specific Methods for Field Data Access --

	SetItems(me : mutable; aItems : mutable HArray1OfAutoDesignGeneralOrgItem);
	Items (me) returns mutable HArray1OfAutoDesignGeneralOrgItem;
	ItemsValue (me; num : Integer) returns AutoDesignGeneralOrgItem;
	NbItems (me) returns Integer;

fields

	items : HArray1OfAutoDesignGeneralOrgItem from StepAP214; -- a SelectType

end AutoDesignApprovalAssignment;
