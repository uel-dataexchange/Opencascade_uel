-- File:	PXCAFDoc_DimTolTool.cdl
-- Created:	Wed Dec 10 12:24:08 2008
-- Author:	Pavel TELKOV
--		<ptv@valenox>
---Copyright:	 Open CASCADE 2008

class DimTolTool from PXCAFDoc inherits Attribute from PDF

is
    Create returns DimTolTool from PXCAFDoc;

end DimTolTool;
