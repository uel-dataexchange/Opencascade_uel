-- File:	BRepFeat_MakePrism.cdl
-- Created:	Tue Feb 13 14:24:53 1996
-- Author:	Jacques GOUSSARD
--		<jag@bravox>
---Copyright:	 Matra Datavision 1996


class MakePrism from BRepFeat inherits Form from BRepFeat

	---Purpose: Describes functions to build prism features.
    	-- These can be depressions or protrusions.
    	-- The semantics of prism feature creation is
    	-- based on the construction of shapes:
    	-- -   along a length
    	-- -   up to a limiting face
    	-- -   from a limiting face to a height.
    	-- The shape defining construction of the prism feature can be 
    	-- either the supporting edge or the concerned area of a face.
    	-- In case of the supporting edge, this contour
    	-- can be attached to a face of the basis shape by
    	-- binding. When the contour is bound to this face,
    	-- the information that the contour will slide on the
    	-- face becomes available to the relevant class methods.
    	-- In case of the concerned area of a face, you
    	-- could, for example, cut it out and move it to a
    	-- different height which will define the limiting
    	-- face of a protrusion or depression.

uses Shape                     from TopoDS,
     Face                      from TopoDS,
     Edge                      from TopoDS,
     DataMapOfShapeListOfShape from TopTools,
     Dir                       from gp,
     DataMapOfShapeShape       from TopTools,
     SequenceOfCurve           from TColGeom,
     Curve                     from Geom,
     StatusError               from BRepFeat
     
raises ConstructionError from Standard

is


    Create

    	returns MakePrism from BRepFeat;
	---Purpose: Builds a prism by projecting a
    	-- wire along the face of a shape. Initializes the prism class.
	---C++: inline


    Create(Sbase     : Shape from TopoDS;
           Pbase     : Shape from TopoDS;
           Skface    : Face  from TopoDS;
	   Direction : Dir   from gp;
           Fuse      : Integer from Standard;
           Modify    : Boolean from Standard)
    
	---Purpose: Builds a prism by projecting a
    	-- wire along the face of a shape. a face Pbase is selected in
    	--   the shape Sbase to serve as the basis for
    	--   the prism. The orientation of the prism will
    	--   be defined by the vector Direction.
    	-- Fuse offers a choice between:
    	-- -   removing matter with a Boolean cut using the setting 0
    	-- -   adding matter with Boolean fusion using the setting 1.
    	--   The sketch face Skface serves to determine
    	-- the type of operation. If it is inside the basis
    	-- shape, a local operation such as glueing can be performed.
    	-- Exceptions
    	-- Standard_ConstructionError if the face
    	-- does not belong to the basis or the prism shape.
    		---C++: inline
    	    	returns MakePrism from BRepFeat;


    Init(me: in out; Sbase     : Shape from TopoDS;
                     Pbase     : Shape from TopoDS;
                     Skface    : Face  from TopoDS;
	             Direction : Dir   from gp;
                     Fuse      : Integer from Standard;
                     Modify    : Boolean from Standard)
    
    	is static;
    	---Purpose: Initializes this algorithm for building prisms along surfaces.
    	-- A face Pbase is selected in the shape Sbase
    	-- to serve as the basis for the prism. The
    	-- orientation of the prism will be defined by the vector Direction.
    	-- Fuse offers a choice between:
    	-- -   removing matter with a Boolean cut using the setting 0
    	-- -   adding matter with Boolean fusion using the setting 1.
    	-- The sketch face Skface serves to determine
    	-- the type of operation. If it is inside the basis
    	-- shape, a local operation such as glueing can be performed.

    Add(me: in out; E: Edge from TopoDS; OnFace: Face from TopoDS)

	---Purpose: Indicates that the edge <E> will slide on the face
	--  <OnFace>. Raises ConstructionError if the  face does not belong to the
	-- basis shape, or the edge to the prismed shape.
    	raises ConstructionError from Standard
	
	is static;


    Perform(me: in out; Length: Real from Standard)
    
    	is static;


    Perform(me: in out; Until:  Shape from TopoDS)
    
    	is static;


    Perform(me: in out; From :  Shape from TopoDS;
                        Until:  Shape from TopoDS)
    
    	is static;
    	---Purpose: Assigns one of the following semantics
    	-- -   to a height Length
    	-- -   to a face Until
    	-- -   from a face From to a height Until.
    	-- Reconstructs the feature topologically according to the semantic option chosen.

    PerformUntilEnd(me: in out)
    
    	is static;
    	--- Purpose: Realizes a semi-infinite prism, limited by the
    	-- position of the prism base. All other faces extend infinitely.

    PerformFromEnd(me: in out; FUntil: Shape from TopoDS)
    
    	is static;
    	---Purpose: Realizes a semi-infinite prism, limited by the face Funtil.


    PerformThruAll(me: in out)
    
    	is static;
    	---Purpose: Builds an infinite prism. The infinite descendants will not be kept in the result.
        
    PerformUntilHeight(me: in out; Until :  Shape from TopoDS;
                        Length:  Real  from Standard)
    
    	is static;
    	---Purpose: Assigns both a limiting shape, Until from
    	-- TopoDS_Shape, and a height, Length at which to stop generation of the prism feature.
        
    Curves(me: in out; S : in out SequenceOfCurve from TColGeom);
    	--- Purpose: Returns the list of curves S parallel to the axis of the prism.   

    BarycCurve(me: in out)    
    	returns Curve from Geom;
    	---Purpose: Generates a curve along the center of mass of the primitive.
fields

    myPbase  : Shape                     from TopoDS;
    mySlface : DataMapOfShapeListOfShape from TopTools;
    myDir    : Dir                       from gp;
    myCurves : SequenceOfCurve           from TColGeom;
    myBCurve : Curve                     from Geom;
    myStatusError : StatusError          from BRepFeat;

end MakePrism;
