-- File:	RWStepRepr_RWExtension.cdl
-- Created:	Wed Jun  4 14:17:23 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWExtension from RWStepRepr

    ---Purpose: Read & Write tool for Extension

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    Extension from StepRepr

is
    Create returns RWExtension from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : Extension from StepRepr);
	---Purpose: Reads Extension

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: Extension from StepRepr);
	---Purpose: Writes Extension

    Share (me; ent : Extension from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWExtension;
