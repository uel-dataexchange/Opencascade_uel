-- File:        BoundaryCurve.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWBoundaryCurve from RWStepGeom

	---Purpose : Read & Write Module for BoundaryCurve

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     BoundaryCurve from StepGeom,
     EntityIterator from Interface

is

	Create returns RWBoundaryCurve;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable BoundaryCurve from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : BoundaryCurve from StepGeom);

	Share(me; ent : BoundaryCurve from StepGeom; iter : in out EntityIterator);

end RWBoundaryCurve;
