-- File:	FuncExtPS.cdl
-- Created:	Wed Jul 24 14:31:49 1991
-- Author:	Michel CHAUVAT
--		<mca@topsn3>
---Copyright:	 Matra Datavision 1991

-- Modified by skv - Thu Sep 30 15:19:59 2004 OCC593


private class FuncExtPS from Extrema

 inherits FunctionSetWithDerivatives from math
    ---Purpose: Fonction permettant de rechercher les extrema de la 
    --          distance entre un point et une surface.

uses    POnSurf           from Extrema,
	SequenceOfPOnSurf from Extrema,
	SequenceOfReal    from TColStd,
	Pnt               from gp,
	Vector            from math,
	Matrix            from math,
	Surface           from Adaptor3d,
    	SurfacePtr        from Adaptor3d

raises  OutOfRange from Standard

is
    Create returns FuncExtPS;

    Create (P: Pnt; S: Surface from Adaptor3d) returns FuncExtPS;
    	---Purpose:

    Initialize(me: in out; S: Surface from Adaptor3d)
    	---Purpose: sets the field mysurf of the function.
    is static;
    
    SetPoint(me: in out; P: Pnt)
    	---Purpose: sets the field mysurf of the function.
    is static;

    ------------------------------------------------------------
    -- In all next methods, an exception is raised if the fields 
    -- were not initialized.

    NbVariables (me) returns Integer;

    NbEquations (me) returns Integer;

    Value (me: in out; UV: Vector; F: out Vector) returns Boolean;
    	---Purpose: Calcul de Fi(U,V).

    Derivatives (me: in out; UV: Vector; DF: out Matrix)
    	returns Boolean;
    	---Purpose: Calcul de Fi'(U,V).

    Values (me: in out; UV: Vector; F: out Vector; DF: out Matrix)
    	returns Boolean;
    	---Purpose: Calcul de Fi(U,V) et Fi'(U,V).

    GetStateNumber (me: in out) returns Integer
    	---Purpose: Memorise l'extremum trouve.
    	is redefined;

    NbExt (me) returns Integer;
    	---Purpose: Renvoie le nombre d'extrema trouves.

    SquareDistance (me; N: Integer) returns Real
    	---Purpose: Renvoie la valeur de la Nieme distance.
    	raises  OutOfRange;
	    	-- si N < 1 ou N > NbExt(me).

    Point (me; N: Integer) returns POnSurf
    	---Purpose: Renvoie le Nieme extremum.
    	raises  OutOfRange;
	    	-- si N < 1 ou N > NbExt(me).

-- Modified by skv - Thu Sep 30 15:19:59 2004 OCC593 Begin
    HasDegIso(me) returns Boolean from Standard;
-- Modified by skv - Thu Sep 30 15:19:59 2004 OCC593 End

    Bidon(me) returns SurfacePtr from Adaptor3d
    is static private;
 
fields
    myP    : Pnt from gp;
    myS    : SurfacePtr from Adaptor3d;

    myU    : Real;          -- valeur courante de U
    myV    : Real;          -- valeur courante de V
    myPs   : Pnt from gp;   -- point courant

    mySqDist: SequenceOfReal    from TColStd;
    myPoint: SequenceOfPOnSurf from Extrema;
    myPinit: Boolean;
    mySinit: Boolean;
    myUIsoIsDeg: Boolean;
    myVIsoIsDeg: Boolean;

end FuncExtPS;
