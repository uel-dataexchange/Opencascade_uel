-- File:	IGESGeom_ToolFlash.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolFlash  from IGESGeom

    ---Purpose : Tool to work on a Flash. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses Flash from IGESGeom,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolFlash;
    ---Purpose : Returns a ToolFlash, ready to work


    ReadOwnParams (me; ent : mutable Flash;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : Flash;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : Flash;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a Flash <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable Flash) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a Flash
    --           (LineFont in Directory Entry forced to Rank = 1)

    DirChecker (me; ent : Flash) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : Flash;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : Flash; entto : mutable Flash;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : Flash;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolFlash;
