-- File:	IntConicQuad.cdl
-- Created:	Thu Aug  6 10:51:07 1992
-- Author:	Laurent BUCHARD
--		<lbr@sdsun2>
---Copyright:	 Matra Datavision 1992


class IntConicQuad from IntAna 

	---Purpose: This class provides the analytic intersection between
	--          a conic defined as an element of gp (Lin,Circ,Elips,
	--          Parab,Hypr) and a quadric as defined in the class
	--          Quadric from IntAna.
	--          The intersection between a conic and a plane is treated
	--          as a special case.
	--          
	--          The result of the intersection are points (Pnt from
	--          gp), associated with the parameter on the conic.
	--          
    	--          A call to an Intersection  L:Lin from gp and 
    	--          SPH: Sphere from gp can be written either : 
    	--               IntAna_IntConicQuad Inter(L,IntAna_Quadric(SPH))
    	--           or :
    	--               IntAna_IntConicQuad Inter(L,SPH) (it is necessary
    	--                  to include IntAna_Quadric.hxx in this case)



uses Pnt     from gp,
     Lin     from gp,
     Circ    from gp,
     Elips   from gp,
     Parab   from gp,
     Hypr    from gp,
     Pln     from gp,
     Quadric from IntAna
     
     

raises NotDone     from StdFail,
       OutOfRange  from Standard,
       DomainError from Standard

is


    Create
    
    	---Purpose: Empty constructor.
    	--          
    
	returns IntConicQuad from IntAna;



    Create(L: Lin from gp; Q: Quadric from IntAna)
    
    	---Purpose: Creates the intersection between a line and a quadric.

    	returns IntConicQuad from IntAna;


    Perform(me:in out; L: Lin from gp; Q: Quadric from IntAna)
    
    	---Purpose: Intersects a line and a quadric.

    	is static;


    Create(C: Circ from gp; Q: Quadric from IntAna)
    
    	---Purpose: Creates the intersection between a circle and a quadric.

    	returns IntConicQuad from IntAna;


    Perform(me: in out; C: Circ from gp; Q: Quadric from IntAna)
    
    	---Purpose: Intersects a circle and a quadric.

    	is static;


    Create(E: Elips from gp; Q: Quadric from IntAna)
    
    	---Purpose: Creates the intersection between an ellipse and a quadric.

    	returns IntConicQuad from IntAna;


    Perform(me:in out; E: Elips from gp; Q: Quadric from IntAna)
    
    	---Purpose: Intersects an ellipse and a quadric.

    	is static;


    Create(P: Parab from gp; Q: Quadric from IntAna)
    
    	---Purpose: Creates the intersection between a parabola and a quadric.

    	returns IntConicQuad from IntAna;


    Perform(me:in out; P: Parab from gp; Q: Quadric from IntAna)
    
    	---Purpose: Intersects a parabola and a quadric.

        is static;


    Create(H: Hypr from gp; Q: Quadric from IntAna)
    
    	---Purpose: Creates the intersection between an hyperbola and
    	--          a quadric.

    	returns IntConicQuad from IntAna;


    Perform(me:in out; H: Hypr from gp; Q: Quadric from IntAna)
    
    	---Purpose: Intersects an hyperbola and a quadric.

    	is static;

----------------------------------------------------------------------
--  Intersection between a Conic from gp and a Pln from IntAna
--  The intersection is computed with Tolerances.
----------------------------------------------------------------------

    Create(L : Lin from gp; P: Pln from gp; 
           Tolang: Real from Standard)
    
	---Purpose: Intersection between a line and a plane.
	--          Tolang is used to determine if the angle between two
	--          vectors is null.
    
    	returns IntConicQuad from IntAna;
	

    Perform(me: in out;
            L : Lin from gp; P: Pln from gp; Tolang: Real from Standard)
    
	---Purpose: Intersects a line and a plane.
	--          Tolang is used to determine if the angle between two
	--          vectors is null.
    
    	is static;
	

    Create(C : Circ from gp; P: Pln from gp; 
           Tolang,Tol: Real from Standard)
    
	---Purpose: Intersection between a circle and a plane.
	--          Tolang is used to determine if the angle between two
	--          vectors is null.
	--          Tol is used to determine if a distance is null.
    
    	returns IntConicQuad from IntAna;


    Perform(me: in out;
            C : Circ from gp; P: Pln from gp; Tolang,Tol: Real from Standard)
    
	---Purpose: Intersects a circle and a plane.
	--          Tolang is used to determine if the angle between two
	--          vectors is null.
	--          Tol is used to determine if a distance is null.
    
    	is static;


    Create(E : Elips from gp; P: Pln from gp; 
           Tolang,Tol: Real from Standard)
    
	---Purpose: Intersection between an ellipse and a plane.
	--          Tolang is used to determine if the angle between two
	--          vectors is null.
	--          Tol is used to determine if a distance is null.
    
    	returns IntConicQuad from IntAna;


    Perform(me: in out;
            E : Elips from gp; P: Pln from gp; Tolang,Tol: Real from Standard)
    
	---Purpose: Intersects an ellipse and a plane.
	--          Tolang is used to determine if the angle between two
	--          vectors is null.
	--          Tol is used to determine if a distance is null.
    
    	is static;


    Create(Pb: Parab from gp; P: Pln from gp; 
           Tolang: Real from Standard)
    
	---Purpose: Intersection between a parabola and a plane.
	--          Tolang is used to determine if the angle between two
	--          vectors is null.
    
    	returns IntConicQuad from IntAna;


    Perform(me: in out;
            Pb: Parab from gp; P: Pln from gp; Tolang: Real from Standard)
    
	---Purpose: Intersects a parabola and a plane.
	--          Tolang is used to determine if the angle between two
	--          vectors is null.
    
    	is static;


    Create(H : Hypr from gp; P: Pln from gp; 
           Tolang: Real from Standard)
    
	---Purpose: Intersection between an hyperbola and a plane.
	--          Tolang is used to determine if the angle between two
	--          vectors is null.
    
    	returns IntConicQuad from IntAna;


    Perform(me: in out;
            H : Hypr from gp; P: Pln from gp; Tolang: Real from Standard)
    
	---Purpose: Intersects an hyperbola and a plane.
	--          Tolang is used to determine if the angle between two
	--          vectors is null.
    
    	is static;


    IsDone(me)
    
    	---Purpose: Returns TRUE if the creation completed.
    	--          
	---C++: inline

    	returns Boolean from Standard
    	is static;


    IsInQuadric(me)
    
    	---Purpose: Returns TRUE if the conic is in the quadric.
    	--          
	---C++: inline

    	returns Boolean from Standard

    	raises NotDone from StdFail
    	--     The exception NotDone is raised if IsDone returns False.
	
	is static;


    IsParallel(me)
    
    	---Purpose: Returns TRUE if the line is in a quadric which
    	--          is parallel to the quadric.
	---C++: inline

    	returns Boolean from Standard

    	raises NotDone from StdFail
    	--     The exception NotDone is raised if IsDone returns False.
	
	is static;


    NbPoints(me)
    
    	---Purpose: Returns the number of intersection point.
    	--          
	---C++: inline

    	returns Integer from Standard

    	raises NotDone      from StdFail, 
               DomainError  from Standard
    	--     The exception NotDone is raised if IsDone returns False.
    	--     The exception DomainError is raised if IsInQuadric returns
    	--          True or IsParallel returns True.

	
	is static;


    Point(me; N: Integer from Standard)
    
    	---Purpose: Returns the point of range N.
    	--          
	---C++: inline
	---C++: return const&

    	returns Pnt from gp

    	raises NotDone     from StdFail, 
               DomainError from Standard, 
               OutOfRange  from Standard
    	--     The exception NotDone is raised if IsDone returns False.
    	--     The exception DomainError is raised if IsInQuadric returns
    	--          True or IsParallel returns true.
    	--     The exception OutOfRange is raised if N<=0 or N>NbPoints.
	
	is static;


    ParamOnConic(me; N: Integer from Standard)
    
    	---Purpose: Returns the parameter on the line of the intersection
    	--          point of range N.
    	--          
	---C++: inline

    	returns Real from Standard
	
	raises NotDone     from StdFail,
               DomainError from Standard,
	       OutOfRange  from Standard
    	--     The exception NotDone is raised if IsDone returns False.
    	--     The exception DomainError is raised if IsInQuadric returns
    	--          True or IsParallel returns true.
    	--     The exception OutOfRange is raised if N<=0 or N>NbPoints.
	
	is static;



fields

    done          : Boolean from Standard;
    parallel      : Boolean from Standard;
    inquadric     : Boolean from Standard;
    
    nbpts         : Integer from Standard;
    
    pnts          : Pnt     from gp [4];
    paramonc      : Real    from Standard [4];

end IntConicQuad;


