-- File:	RWStepShape_RWConnectedFaceSubSet.cdl
-- Created:	Fri Jan  4 17:42:43 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWConnectedFaceSubSet from RWStepShape

    ---Purpose: Read & Write tool for ConnectedFaceSubSet

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ConnectedFaceSubSet from StepShape

is
    Create returns RWConnectedFaceSubSet from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ConnectedFaceSubSet from StepShape);
	---Purpose: Reads ConnectedFaceSubSet

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ConnectedFaceSubSet from StepShape);
	---Purpose: Writes ConnectedFaceSubSet

    Share (me; ent : ConnectedFaceSubSet from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWConnectedFaceSubSet;
