-- File:	GeomLib_IsPlanarSurface.cdl
-- Created:	Mon Nov 23 11:01:50 1998
-- Author:	Philippe MANGIN
--		<pmn@sgi29>
---Copyright:	 Matra Datavision 1998


class IsPlanarSurface from GeomLib 

	---Purpose: Find if a surface is a planar  surface.          

uses 
  Surface  from  Geom, 
  Pln     from  gp

raises 
  NotDone  from  StdFail

is 
  Create(S  :  Surface;  Tol  :  Real  =  1.0e-7) 
  returns  IsPlanarSurface  from  GeomLib; 
   
  IsPlanar(me)  
  ---Purpose: Return if the Surface is a plan
  returns  Boolean; 
   
  Plan(me)   
  ---Purpose: Return the plan definition        
  ---C++: return const &     
  returns  Pln  from  gp 
  raises  NotDone;  --  if  <me>  is  not  Planar

fields 
  myPlan  :  Pln  from  gp; 
  IsPlan  :  Boolean;

end IsPlanarSurface;
