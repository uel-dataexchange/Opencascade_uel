-- File:	PTopoDS_Solid.cdl
-- Created:	Wed May  5 16:57:09 1993
-- Author:	Remi LEQUETTE
--		<rle@sdsun1>
---Copyright:	 Matra Datavision 1993



class Solid from PTopoDS inherits HShape from PTopoDS

is
    Create returns mutable Solid from PTopoDS;
    ---Level: Internal 

end Solid;
