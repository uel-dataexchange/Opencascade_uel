-- File:	StepFEA_ParametricCurve3dElementCoordinateSystem.cdl
-- Created:	Thu Dec 12 17:51:07 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class ParametricCurve3dElementCoordinateSystem from StepFEA
inherits FeaRepresentationItem from StepFEA

    ---Purpose: Representation of STEP entity ParametricCurve3dElementCoordinateSystem

uses
    HAsciiString from TCollection,
    ParametricCurve3dElementCoordinateDirection from StepFEA

is
    Create returns ParametricCurve3dElementCoordinateSystem from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aDirection: ParametricCurve3dElementCoordinateDirection from StepFEA);
	---Purpose: Initialize all fields (own and inherited)

    Direction (me) returns ParametricCurve3dElementCoordinateDirection from StepFEA;
	---Purpose: Returns field Direction
    SetDirection (me: mutable; Direction: ParametricCurve3dElementCoordinateDirection from StepFEA);
	---Purpose: Set field Direction

fields
    theDirection: ParametricCurve3dElementCoordinateDirection from StepFEA;

end ParametricCurve3dElementCoordinateSystem;
