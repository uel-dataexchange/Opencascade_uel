-- File:	StepSelect_StepType.cdl
-- Created:	Thu Dec 22 09:38:35 1994
-- Author:	Christian CAILLET
--		<cky@anion>
---Copyright:	 Matra Datavision 1994


class StepType  from StepSelect    inherits Signature  from IFSelect

    ---Purpose : StepType is a Signature specific to Step definitions : it
    --           considers the type as defined in STEP Schemas, the same which
    --           is used in files.
    --           For a Complex Type, if its definition is known, StepType
    --           produces the list of basic types, separated by commas, the
    --           whole between brackets : "(TYPE1,TYPE2..)".
    --           If its precise definition is not known (simply it is known as
    --           Complex, it can be recognised, but the list is produced at
    --           Write time only), StepType produces : "(..COMPLEX TYPE..)"

uses CString, Transient, AsciiString from TCollection,
     Protocol from Interface, InterfaceModel,
     Protocol from StepData,  WriterLib from StepData

raises InterfaceError

is

    Create returns mutable StepType;
    ---Purpose : Creates a Signature for Step Type. Protocol is undefined here,
    --           hence no Signature may yet be produced. The StepType signature
    --           requires a Protocol before working

    SetProtocol (me : mutable; proto : Protocol from Interface)
    ---Purpose : Sets the StepType signature to work with a Protocol : this
    --           initialises the library
    	raises InterfaceError;
    --           Error if the Protocol is not from StepData

    Value (me; ent : any Transient; model : InterfaceModel) returns CString;
    ---Purpose : Returns the Step Type defined from the Protocol (see above).
    --           If <ent> is not recognised, produces "..NOT FROM SCHEMA <name>.."

fields

    theproto : Protocol  from StepData;
    thelib   : WriterLib from StepData is protected;

end StepType;
