-- File:	PDataStd_Placement.cdl
-- Created:	Tue Jul 29 13:49:37 1997
-- Author:	Denis PASCAL 
-- modified     Sergey Zaritchny
---Copyright:	 Matra Datavision 1997


class Placement from PDataXtd inherits Attribute from PDF

	---Purpose: 

    
is

    Create returns mutable Placement from  PDataXtd;
    

end Placement;
