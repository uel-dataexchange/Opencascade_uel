-- File:	TNaming_UsedShapes.cdl
-- Created:	Wed Feb  5 09:55:14 1997
-- Author:	Yves FRICAUD
--		<yfr@claquox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


private class UsedShapes from TNaming inherits Attribute from TDF

	---Purpose: Set of Shapes Used in a Data from TDF
	--          Only one instance by Data, it always
	--          Stored as Attribute of The Root.

uses
    GUID                      from Standard,
    DataMapOfShapePtrRefShape from TNaming,
    RelocationTable           from TDF,
    AttributeIndexedMap       from TDF,
    Attribute                 from TDF,
    AttributeDelta            from TDF, 
    DeltaOnAddition           from TDF, 
    DeltaOnRemoval            from TDF,
    Delta                     from TDF,
    DataSet	              from TDF

is

    Create returns mutable UsedShapes from TNaming 
    is private;

    Destroy(me : mutable);
    ---C++: alias ~

    Map (me: mutable) returns DataMapOfShapePtrRefShape from TNaming;
    	---C++: return &
    	---C++: inline

    ID(me) returns GUID from Standard
    is redefined static;
	---Purpose: Returns the ID of the attribute.
	---C++: inline 	
	---C++: return const &             	
  
    GetID(myclass) returns GUID from Standard;
	---Purpose: Returns the ID: 2a96b614-ec8b-11d0-bee7-080009dc3333.
    	---C++: return const &
    
    BackupCopy(me) returns mutable Attribute from TDF
    is redefined;
	---Purpose: Copies  the attribute  contents into  a  new other
	--          attribute. It is used by Backup().

    Restore(me: mutable; anAttribute : Attribute from TDF)
    is redefined;
	---Purpose: Restores the contents from <anAttribute> into this
	--          one. It is used when aborting a transaction.

    BeforeRemoval(me: mutable)
    	is redefined;
	---Purpose: Clears the table.

    AfterUndo(me: mutable;
    	      anAttDelta : AttributeDelta from TDF;
    	      forceIt : Boolean from Standard = Standard_False)
    	returns Boolean from Standard
    	is redefined;
	---Purpose: Something to do after applying <anAttDelta>.

 
    ---Category: Delta generation
    --           =================================================

    DeltaOnAddition(me)
    	returns DeltaOnAddition from TDF is redefined;
    	---Purpose : this method returns a null handle (no delta).
    	


    DeltaOnRemoval(me)
    	returns DeltaOnRemoval from TDF is redefined;
    	---Purpose : this method returns a null handle (no delta).
    	


    -- Copy use methods
    -- ----------------

    NewEmpty(me)
    	returns mutable Attribute from TDF
    	is redefined;
	---Purpose: Returns an new empty attribute from the good end
	--          type. It is used by the copy algorithm.

    Paste(me;
    	  intoAttribute    : mutable Attribute from TDF;
	  aRelocTationable : mutable RelocationTable from TDF)
 	is redefined;
	---Purpose: This method is different from the "Copy" one,
	--          because it is used when copying an attribute from
	--          a source structure into a target structure. This
	--          method pastes the current attribute to the label
	--          corresponding to the insertor. The pasted
	--          attribute may be a brand new one or a new version
	--          of the previous one.
 
    References(me; aDataSet : DataSet from TDF)
    	is redefined;
	---Purpose: Adds the directly referenced attributes and labels
	--          to <aDataSet>. "Directly" means we have only to
	--          look at the first level of references.
	--          
	--          For this, use only the AddLabel() & AddAttribute()
	--          from DataSet and do not try to modify information
	--          previously stored in <aDataSet>.


    -- Miscelleaneous
    -- --------------
    Dump(me; anOS : in out OStream from Standard)
    	returns OStream from Standard
    	is redefined ;
	---Purpose: Dumps the attribute on <aStream>.
    	---C++ : return &


fields
    myMap : DataMapOfShapePtrRefShape from TNaming;
    
friends
    class Builder from TNaming

end UsedShapes;
