-- File:	TopoDSToStep_MakeGeometricCurveSet.cdl
-- Created:	Fri Mar 17 10:54:55 1995
-- Author:	Dieter THIEMANN
--		<dth@cinox>
---Copyright:	 Matra Datavision 1995


class MakeGeometricCurveSet from TopoDSToStep inherits
    Root from TopoDSToStep

    ---Purpose: This class implements the mapping between a Shape 
    --          from TopoDS and a GeometricCurveSet from StepShape in order
    --          to create a GeometricallyBoundedWireframeRepresentation.
  
uses Shape from TopoDS,
     GeometricCurveSet from StepShape,
     FinderProcess from Transfer
          
raises NotDone from StdFail
     
is 

Create ( SH : Shape from TopoDS;
         FP : mutable FinderProcess from Transfer)
        returns MakeGeometricCurveSet;

Value (me) returns GeometricCurveSet from StepShape
    raises NotDone
    is static;
    ---C++: return const&

fields

    theGeometricCurveSet : GeometricCurveSet from StepShape;
    
    
end MakeGeometricCurveSet;    
