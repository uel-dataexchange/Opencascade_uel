-- File:	PGeom_BezierCurve.cdl
-- Created:	Mon Feb 22 18:59:59 1993
-- Author:	Philippe DAUTRY
--		<fid@phobox>
-- Copyright:	 Matra Datavision 1993


class BezierCurve from PGeom inherits BoundedCurve from PGeom

        ---Purpose : Defines a rational or non rational Bezier curve.
        --         
	---See Also : BezierCurve from Geom.

uses  HArray1OfReal from PColStd,
      HArray1OfPnt  from PColgp

is 


  Create returns mutable BezierCurve from PGeom;
        ---Purpose : Creates a non rational  Bezier curve with default
        --         values.
    	---Level: Internal 

  Create(aPoles    : HArray1OfPnt;
         aWeights  : HArray1OfReal;
	 aRational : Boolean from Standard)
     returns mutable BezierCurve from PGeom;
        ---Purpose : Creates a non rational Bezier curve with a set of
        --         poles aCurvePoles and a set of weights aPoleWeight.
    	---Level: Internal 


  Rational (me: mutable; aRational: Boolean from Standard);
        ---Purpose : Set the value of the field rational with <aRational>.
    	---Level: Internal 


  Rational (me) returns Boolean;
        ---Purpose : Returns the value of the field rational.
    	---Level: Internal 


  Poles (me: mutable; aPoles : HArray1OfPnt from PColgp);
        ---Purpose : Set the value of the field poles with <aPoles>.
    	---Level: Internal 


  Poles (me) returns HArray1OfPnt from PColgp;
        ---Purpose : Returns the value of the field poles.
    	---Level: Internal 


  Weights (me: mutable; aWeights : HArray1OfReal from PColStd);
        ---Purpose : Set the value of the field weights.
    	---Level: Internal 


  Weights (me)returns HArray1OfReal from PColStd;
        ---Purpose : Returns the value of the field weights.
    	---Level: Internal 


fields

   rational : Boolean from Standard;
   poles    : HArray1OfPnt  from PColgp;
   weights  : HArray1OfReal from PColStd;

end;
