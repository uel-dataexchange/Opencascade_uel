-- File:	StepElement_MeasureOrUnspecifiedValueMember.cdl
-- Created:	Tue Dec 10 18:12:58 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V2.0
-- Copyright:	Open CASCADE 2002

class MeasureOrUnspecifiedValueMember from StepElement
inherits SelectNamed from StepData

    ---Purpose: Representation of member for  STEP SELECT type MeasureOrUnspecifiedValue

is
    Create returns MeasureOrUnspecifiedValueMember from StepElement;
	---Purpose: Empty constructor

    HasName (me) returns Boolean  is redefined;
	---Purpose: Returns True if has name

    Name (me) returns CString  is redefined;
	---Purpose: Returns set name 

    SetName (me : mutable; name : CString)  returns Boolean  is redefined;
	---Purpose: Set name 

    Matches (me; name : CString) returns Boolean  is redefined;
	---Purpose : Tells if the name of a SelectMember matches a given one;

fields

    mycase : Integer;

end MeasureOrUnspecifiedValueMember;
