-- File:        PresentationSet.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPresentationSet from RWStepVisual

	---Purpose : Read & Write Module for PresentationSet

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PresentationSet from StepVisual

is

	Create returns RWPresentationSet;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PresentationSet from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : PresentationSet from StepVisual);

end RWPresentationSet;
