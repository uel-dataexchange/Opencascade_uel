-- File:	StepDimTol_PerpendicularityTolerance.cdl
-- Created:	Wed Jun  4 13:34:34 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class PerpendicularityTolerance from StepDimTol
inherits GeometricToleranceWithDatumReference from StepDimTol

    ---Purpose: Representation of STEP entity PerpendicularityTolerance

uses
    HAsciiString from TCollection,
    MeasureWithUnit from StepBasic,
    ShapeAspect from StepRepr,
    HArray1OfDatumReference from StepDimTol

is
    Create returns PerpendicularityTolerance from StepDimTol;
	---Purpose: Empty constructor

end PerpendicularityTolerance;
