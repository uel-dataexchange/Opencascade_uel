-- File:	RWStepDimTol_RWPerpendicularityTolerance.cdl
-- Created:	Wed Jun  4 13:34:34 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWPerpendicularityTolerance from RWStepDimTol

    ---Purpose: Read & Write tool for PerpendicularityTolerance

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    PerpendicularityTolerance from StepDimTol

is
    Create returns RWPerpendicularityTolerance from RWStepDimTol;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : PerpendicularityTolerance from StepDimTol);
	---Purpose: Reads PerpendicularityTolerance

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: PerpendicularityTolerance from StepDimTol);
	---Purpose: Writes PerpendicularityTolerance

    Share (me; ent : PerpendicularityTolerance from StepDimTol;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWPerpendicularityTolerance;
