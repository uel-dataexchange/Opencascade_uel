-- File:	StepFEA_CurveElementEndRelease.cdl
-- Created:	Thu Dec 12 17:51:04 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class CurveElementEndRelease from StepFEA
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity CurveElementEndRelease

uses
    CurveElementEndCoordinateSystem from StepFEA,
    HArray1OfCurveElementEndReleasePacket from StepElement

is
    Create returns CurveElementEndRelease from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aCoordinateSystem: CurveElementEndCoordinateSystem from StepFEA;
                       aReleases: HArray1OfCurveElementEndReleasePacket from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    CoordinateSystem (me) returns CurveElementEndCoordinateSystem from StepFEA;
	---Purpose: Returns field CoordinateSystem
    SetCoordinateSystem (me: mutable; CoordinateSystem: CurveElementEndCoordinateSystem from StepFEA);
	---Purpose: Set field CoordinateSystem

    Releases (me) returns HArray1OfCurveElementEndReleasePacket from StepElement;
	---Purpose: Returns field Releases
    SetReleases (me: mutable; Releases: HArray1OfCurveElementEndReleasePacket from StepElement);
	---Purpose: Set field Releases

fields
    theCoordinateSystem: CurveElementEndCoordinateSystem from StepFEA;
    theReleases: HArray1OfCurveElementEndReleasePacket from StepElement;

end CurveElementEndRelease;
