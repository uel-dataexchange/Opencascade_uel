-- File:        Conic.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWConic from RWStepGeom

	---Purpose : Read & Write Module for Conic

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Conic from StepGeom,
     EntityIterator from Interface

is

	Create returns RWConic;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Conic from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : Conic from StepGeom);

	Share(me; ent : Conic from StepGeom; iter : in out EntityIterator);

end RWConic;
