-- File:        PolyLoop.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPolyLoop from RWStepShape

	---Purpose : Read & Write Module for PolyLoop

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PolyLoop from StepShape,
     EntityIterator from Interface

is

	Create returns RWPolyLoop;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PolyLoop from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : PolyLoop from StepShape);

	Share(me; ent : PolyLoop from StepShape; iter : in out EntityIterator);

end RWPolyLoop;
