-- File:        PresentationRepresentation.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPresentationRepresentation from RWStepVisual

	---Purpose : Read & Write Module for PresentationRepresentation

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PresentationRepresentation from StepVisual,
     EntityIterator from Interface

is

	Create returns RWPresentationRepresentation;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PresentationRepresentation from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : PresentationRepresentation from StepVisual);

	Share(me; ent : PresentationRepresentation from StepVisual; iter : in out EntityIterator);

end RWPresentationRepresentation;
