-- File:	StepDimTol_GeometricTolerance.cdl
-- Created:	Wed Jun  4 13:34:35 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class GeometricTolerance from StepDimTol
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity GeometricTolerance

uses
    HAsciiString from TCollection,
    MeasureWithUnit from StepBasic,
    ShapeAspect from StepRepr

is
    Create returns GeometricTolerance from StepDimTol;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       aDescription: HAsciiString from TCollection;
                       aMagnitude: MeasureWithUnit from StepBasic;
                       aTolerancedShapeAspect: ShapeAspect from StepRepr);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

    Magnitude (me) returns MeasureWithUnit from StepBasic;
	---Purpose: Returns field Magnitude
    SetMagnitude (me: mutable; Magnitude: MeasureWithUnit from StepBasic);
	---Purpose: Set field Magnitude

    TolerancedShapeAspect (me) returns ShapeAspect from StepRepr;
	---Purpose: Returns field TolerancedShapeAspect
    SetTolerancedShapeAspect (me: mutable; TolerancedShapeAspect: ShapeAspect from StepRepr);
	---Purpose: Set field TolerancedShapeAspect

fields
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection;
    theMagnitude: MeasureWithUnit from StepBasic;
    theTolerancedShapeAspect: ShapeAspect from StepRepr;

end GeometricTolerance;
