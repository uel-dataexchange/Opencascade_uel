-- File:	SelectionIterator.cdl
-- Created:	Tue Nov 17 15:18:39 1992
-- Author:	Christian CAILLET
--		<cky@topsn2>
---Copyright:	 Matra Datavision 1992


class SelectionIterator  from IFSelect

    ---Purpose : Defines an Iterator on a list of Selections

uses Selection, HSeqOfSelection, TSeqOfSelection

raises NoSuchObject

is

    Create  returns SelectionIterator;
    ---Purpose : Creates an empty iterator, ready to be filled

    Create (sel : Selection) returns SelectionIterator;
    ---Purpose : Creates an iterator from a Selection : it lists the Selections
    --           from which <sel> depends (given by its method FillIterator)

    AddFromIter (me : in out;  iter : in out SelectionIterator)  is static;
    ---Purpose : Adds to an iterator the content of another one
    --           (each selection is present only once in the result)

    AddItem     (me : in out; sel : any Selection)               is static;
    ---Purpose : Adds a Selection to an iterator (if not yet noted)

    AddList     (me : in out; list : TSeqOfSelection)            is static;
    ---Purpose : Adds a list of Selections to an iterator (this list comes
    --           from the description of a Selection or a Dispatch, etc...)


    More (me) returns Boolean  is static;
    ---Purpose : Returns True if there are more Selections to get

    Next (me : in out)  is static;
    ---Purpose : Sets iterator to the next item

    Value (me) returns any Selection  raises NoSuchObject  is static;
    ---Purpose : Returns the current Selction beeing iterated
    --           Error if count of Selection has been passed
    ---C++ : return const &

fields

    thecurr : Integer;
    thelist : HSeqOfSelection;

end SelectionIterator;
