-- File:	TDF_DeltaOnResume.cdl
--      	---------------------
-- Author:	DAUTRY Philippe
--		<fid@fox.paris1.matra-dtv.fr>
---Copyright:	 MATRA DATAVISION 1998

---Version:	0.0
---History:	Version	Date		Purpose
--		0.0	Jul  6 1998	Creation
--		1.0	Jul  6 1998	Separation Forget/Resume

class DeltaOnResume from TDF inherits AttributeDelta from TDF

	---Purpose: This class provides default services for an
	--          AttributeDelta on an Resume action.
	--          
	--          Applying this AttributeDelta means FORGETTING its
	--          attribute.

uses

    Attribute from TDF

is

    Create(anAtt : Attribute from TDF)
    	returns mutable DeltaOnResume from TDF;
	---Purpose: Creates a TDF_DeltaOnResume.

    Apply (me : mutable)
    	is redefined static;
    	---Purpose: Applies the delta to the attribute.

end DeltaOnResume;
