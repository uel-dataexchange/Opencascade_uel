-- File:	RWStepDimTol_RWPositionTolerance.cdl
-- Created:	Wed Jun  4 13:34:34 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWPositionTolerance from RWStepDimTol

    ---Purpose: Read & Write tool for PositionTolerance

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    PositionTolerance from StepDimTol

is
    Create returns RWPositionTolerance from RWStepDimTol;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : PositionTolerance from StepDimTol);
	---Purpose: Reads PositionTolerance

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: PositionTolerance from StepDimTol);
	---Purpose: Writes PositionTolerance

    Share (me; ent : PositionTolerance from StepDimTol;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWPositionTolerance;
