-- File:        MDataStd_TickStorageDriver.cdl
-- Created:     May 29 11:40:00 2007
-- Author:      Vlad Romashko
--  	    	<vladislav.romashko@opencascade.com>
-- Copyright:   Open CASCADE

class TickStorageDriver from MDataStd inherits ASDriver from MDF

uses 

    SRelocationTable from MDF,
    Attribute        from TDF,
    Attribute        from PDF, 
    MessageDriver    from CDM

is

    Create (theMessageDriver : MessageDriver from CDM) 
    returns mutable TickStorageDriver from MDataStd;

    VersionNumber(me) 
    returns Integer from Standard;

    SourceType(me) 
    returns Type from Standard;
    ---Purpose: Returns the type Tick from TDataStd.

    NewEmpty(me) 
    returns mutable Attribute from PDF;

    Paste(me;
    	  Source     :         Attribute from TDF;
    	  Target     : mutable Attribute from PDF;
    	  RelocTable : SRelocationTable from MDF);

end TickStorageDriver;

