-- File:	RWStepRepr_RWMaterialDesignation.cdl
-- Created:	Fri Jul 24 15:48:22 1998
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1998


class RWMaterialDesignation from RWStepRepr

	---Purpose : Read & Write Module for MaterialDesignation

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     MaterialDesignation from StepRepr,
     EntityIterator from Interface

is

	Create returns RWMaterialDesignation;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable MaterialDesignation from StepRepr);

	WriteStep (me; SW : in out StepWriter; ent : MaterialDesignation from StepRepr);

	Share(me; ent : MaterialDesignation from StepRepr; iter : in out EntityIterator);

end RWMaterialDesignation;
