-- File:	GeomFill_CurveAndTrihedron.cdl
-- Created:	Tue Dec  2 11:51:44 1997
-- Author:	Philippe MANGIN
--		<pmn@sgi29>
---Copyright:	 Matra Datavision 1997


class CurveAndTrihedron from GeomFill  
inherits  LocationLaw from GeomFill 

	---Purpose: Define location law with an TrihedronLaw and an
	--           curve           
	--        Definition Location is :            
	--         transformed  section   coordinates  in  (Curve(v)),
	--         (Normal(v),   BiNormal(v), Tangente(v))) systeme are
	--         the  same like section  shape coordinates in 
	--         (O,(OX, OY, OZ)) systeme.
	
uses  
 TrihedronLaw   from GeomFill,
 HCurve         from  Adaptor3d,
 Mat            from  gp, 
 Vec            from  gp,  
 Pnt            from  gp,
 Array1OfReal   from TColStd,
 Array1OfPnt2d  from TColgp, 
 Array1OfVec2d  from TColgp, 
 Shape          from GeomAbs 
 
raises  OutOfRange 

is  
  Create(Trihedron  :  TrihedronLaw from GeomFill) 
    returns CurveAndTrihedron from GeomFill; 

  SetCurve(me : mutable;  C  :  HCurve  from  Adaptor3d) 
   is  redefined;     
    
  GetCurve(me)   
   returns HCurve  from  Adaptor3d  
    ---C++: return const &      
   is redefined;  
    
  SetTrsf(me  :  mutable;  Transfo  :  Mat  from  gp) 
   ---Purpose:  Set a transformation Matrix like   the law M(t) become
   --          Mat * M(t)
  is  redefined;
   
  Copy(me)   
    returns  LocationLaw  from  GeomFill          
  is redefined;
   
-- 
--========== To compute Location and derivatives Location
--              
   D0(me : mutable; 
      Param: Real; 
      M    : out  Mat  from  gp; 
      V    : out  Vec  from  gp)
      ---Purpose: compute Location and 2d points        
   returns Boolean  is  redefined;
 

   D0(me : mutable; 
      Param: Real; 
      M    : out  Mat  from  gp; 
      V    : out  Vec  from  gp;
      Poles2d  : out Array1OfPnt2d from TColgp)
      ---Purpose: compute Location and 2d points        
   returns Boolean  is  redefined;
	
   D1(me : mutable;
      Param: Real; 
      M    : out  Mat  from  gp; 
      V    : out  Vec  from  gp; 
      DM   : out  Mat  from  gp; 
      DV   : out  Vec  from  gp;             
      Poles2d  : out Array1OfPnt2d from TColgp;
      DPoles2d : out Array1OfVec2d from TColgp)
      ---Purpose: compute location 2d  points and  associated
      --          first derivatives.         
      --  Warning : It used only for C1 or C2 aproximation
   returns Boolean   
   is  redefined; 
   
   D2(me : mutable;
      Param: Real;
      M    : out  Mat  from  gp; 
      V    : out  Vec  from  gp; 
      DM   : out  Mat  from  gp; 
      DV   : out  Vec  from  gp;   
      D2M  : out  Mat  from  gp; 
      D2V  : out  Vec  from  gp;  
      Poles2d   : out Array1OfPnt2d from TColgp;
      DPoles2d  : out Array1OfVec2d from TColgp;
      D2Poles2d : out Array1OfVec2d from TColgp)      
      ---Purpose: compute location 2d  points and associated
      --          first and seconde  derivatives.
      --  Warning : It used only for C2 aproximation
   returns Boolean
   is  redefined;
           
--
--  =================== Management  of  continuity  ===================
--                 
    NbIntervals(me; S : Shape from GeomAbs) 
	---Purpose: Returns  the number  of  intervals for  continuity
	--          <S>. 
        --          May be one if Continuity(me) >= <S>
   returns Integer  is  redefined;

   Intervals(me; T : in out Array1OfReal from TColStd; 
    	         S : Shape from GeomAbs)
	---Purpose: Stores in <T> the  parameters bounding the intervals
	--          of continuity <S>.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
    raises
    	OutOfRange from Standard 
    is redefined;  
     
    	
   SetInterval(me: mutable; First, Last: Real from Standard)    
	---Purpose: Sets the bounds of the parametric interval on 
	--          the function
	--          This determines the derivatives in these values if the
	--          function is not Cn.
    	is redefined; 
   
    GetInterval(me; First, Last: out  Real from Standard)    
	---Purpose: Gets the bounds of the parametric interval on 
	--          the function
        is redefined;  
	 
    GetDomain(me; First, Last: out  Real from Standard)  
    	---Purpose: Gets the bounds of the function parametric domain.
    	--  Warning: This domain it is  not modified by the
    	--          SetValue method         
        is  redefined;

--  ===================  To help   computation of  Tolerance   ===============
--  
--  Evaluation of error,  in  2d space,  or  on composed function,  is
--  difficult.  The  following methods can  help the  approximation to
--  make good evaluation and use good tolerances.
--      
--      It is not necessary for the following informations to be very
--      precise. A fast evaluation is sufficient.
       
   
  GetMaximalNorm(me  :  mutable)
    ---Purpose:  Get the maximum Norm  of the matrix-location part.  It
    --           is usful to find an good Tolerance to approx M(t).  
  returns Real
  is  redefined;  
   
  GetAverageLaw(me :  mutable;   
                AM: out Mat  from  gp;   
                AV: out Vec  from  gp) 
     ---Purpose: Get average value of M(t) and V(t) it is usfull to 
     --          make fast approximation of rational  surfaces.        
  is  redefined; 
  
-- 
-- To find elementary sweep
-- 
  IsTranslation(me; Error  :  out  Real)  
  ---Purpose: Say if the Location  Law, is an translation of  Location
   -- The default implementation is " returns False ". 
  returns  Boolean
  is redefined;
     
  IsRotation(me; Error  :  out  Real ) 
   ---Purpose: Say if the Location  Law, is a rotation of Location
    -- The default implementation is " returns False ". 
  returns  Boolean 
  is  redefined;  
   
  Rotation(me; Center  :  out  Pnt  from  gp) 
  is redefined;
  
fields 
  WithTrans:  Boolean  from  Standard; 
  myLaw    :  TrihedronLaw  from  GeomFill; 
  myCurve  :  HCurve  from  Adaptor3d;  
  myTrimmed:  HCurve  from  Adaptor3d;  
  Point    :  Pnt  from  gp; 
  V1,  V2,  V3  :  Vec  from  gp;  
  Trans    :  Mat  from gp; 
end CurveAndTrihedron;














