-- File:        CompoundRepresentationItem.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWCompoundRepresentationItem from RWStepRepr

	---Purpose : Read & Write Module for CompoundRepresentationItem

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     EntityIterator from Interface,
     CompoundRepresentationItem from StepRepr

is

	Create returns RWCompoundRepresentationItem;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable CompoundRepresentationItem from StepRepr);

	WriteStep (me; SW : in out StepWriter; ent : CompoundRepresentationItem from StepRepr);

	Share (me; ent : CompoundRepresentationItem from StepRepr;
               iter: in out EntityIterator from Interface);
        ---Purpose: Fills data for graph (shared items)

end RWCompoundRepresentationItem;
