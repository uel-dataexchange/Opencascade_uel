-- File:	IGESAppli_ToolNodalDisplAndRot.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolNodalDisplAndRot  from IGESAppli

    ---Purpose : Tool to work on a NodalDisplAndRot. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses NodalDisplAndRot from IGESAppli,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolNodalDisplAndRot;
    ---Purpose : Returns a ToolNodalDisplAndRot, ready to work


    ReadOwnParams (me; ent : mutable NodalDisplAndRot;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : NodalDisplAndRot;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : NodalDisplAndRot;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a NodalDisplAndRot <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : NodalDisplAndRot) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : NodalDisplAndRot;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : NodalDisplAndRot; entto : mutable NodalDisplAndRot;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : NodalDisplAndRot;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolNodalDisplAndRot;
