-- File:	TopOpeBRepBuild_FaceAreaBuilder.cdl
-- Created:	Thu Dec 21 17:07:40 1995
-- Author:	Jean Yves LEBEY
--		<jyl@meteox>
---Copyright:	 Matra Datavision 1995

class FaceAreaBuilder from TopOpeBRepBuild 
    inherits Area2dBuilder from TopOpeBRepBuild

---Purpose: 
-- The FaceAreaBuilder algorithm is used to construct Faces from a LoopSet,
-- where the Loop is the composite topological object of the boundary,
-- here wire or block of edges.
-- The LoopSet gives an iteration on Loops.
-- For each Loop  it indicates if it is on the boundary (wire) or if it
-- results from  an interference (block of edges).
-- The result of the FaceAreaBuilder is an iteration on areas.
-- An area is described by a set of Loops.

uses

    LoopSet from TopOpeBRepBuild,
    LoopClassifier from TopOpeBRepBuild
    
is

    Create returns FaceAreaBuilder;

    Create(LS : in out LoopSet; LC : in out LoopClassifier;
    	   ForceClass : Boolean = Standard_False) returns FaceAreaBuilder;
    ---Purpose: Creates a FaceAreaBuilder to build faces on
    -- the (wires,blocks of edge) of <LS>, using the classifier <LC>.
    
    InitFaceAreaBuilder(me: in out;
    	    	   	LS : in out LoopSet; LC : in out LoopClassifier;
    	    	    	ForceClass : Boolean = Standard_False) is static;
		    
end FaceAreaBuilder from TopOpeBRepBuild;
