-- File:        TransitionalShapeRepresentation.cdl
-- Created:     Mon Dec  4 12:02:32 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWTransitionalShapeRepresentation from RWStepShape

	---Purpose : Read & Write Module for TransitionalShapeRepresentation

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     TransitionalShapeRepresentation from StepShape,
     EntityIterator from Interface

is

	Create returns RWTransitionalShapeRepresentation;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable TransitionalShapeRepresentation from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : TransitionalShapeRepresentation from StepShape);

	Share(me; ent : TransitionalShapeRepresentation from StepShape; iter : in out EntityIterator);

end RWTransitionalShapeRepresentation;
