-- File:	StepElement_SurfaceElementPurpose.cdl
-- Created:	Tue Dec 10 18:13:04 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V2.0
-- Copyright:	Open CASCADE 2002

class SurfaceElementPurpose from StepElement
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type SurfaceElementPurpose

uses
    SelectMember from StepData,
    EnumeratedSurfaceElementPurpose from StepElement,
    HAsciiString from TCollection

is
    Create returns SurfaceElementPurpose from StepElement;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of SurfaceElementPurpose select type
	--          return 0 

    CaseMem (me; ent: SelectMember from StepData) returns Integer is redefined;
	---Purpose: Recognizes a items of select member SurfaceElementPurposeMember
	--          1 -> EnumeratedSurfaceElementPurpose
	--          2 -> ApplicationDefinedElementPurpose
	--          0 else


     NewMember(me) returns SelectMember from StepData is redefined;
	---Purpose: Returns a new select member the type SurfaceElementPurposeMember

    SetEnumeratedSurfaceElementPurpose(me: in out; aVal :EnumeratedSurfaceElementPurpose from StepElement);
	---Purpose: Set Value for EnumeratedSurfaceElementPurpose

    EnumeratedSurfaceElementPurpose (me) returns EnumeratedSurfaceElementPurpose from StepElement;
	---Purpose: Returns Value as EnumeratedSurfaceElementPurpose (or Null if another type)

    SetApplicationDefinedElementPurpose(me: in out; aVal :HAsciiString from TCollection);
	---Purpose: Set Value for ApplicationDefinedElementPurpose

    ApplicationDefinedElementPurpose (me) returns HAsciiString from TCollection;
	---Purpose: Returns Value as ApplicationDefinedElementPurpose (or Null if another type)

end SurfaceElementPurpose;
