-- File:	TopoDS_Shell.cdl
-- Created:	Mon Dec 17 11:12:03 1990
-- Author:	Remi Lequette
---Copyright:	 Matra Datavision 1990, 1992


class Shell from TopoDS inherits Shape from TopoDS

	---Purpose: Describes a shell which
-- - references an underlying shell with the potential to
--   be given a location and an orientation
-- - has a location for the underlying shell, giving its
--   placement in the local coordinate system
-- - has an orientation for the underlying shell, in terms
--   of its geometry (as opposed to orientation in relation to other shapes).

is
    Create returns Shell from TopoDS;
    ---C++: inline
	---Purpose: Constructs an Undefined Shell.

end Shell;
