-- File:	RWStepBasic_RWGroupAssignment.cdl
-- Created:	Wed May 10 15:09:07 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWGroupAssignment from RWStepBasic

    ---Purpose: Read & Write tool for GroupAssignment

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    GroupAssignment from StepBasic

is
    Create returns RWGroupAssignment from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : GroupAssignment from StepBasic);
	---Purpose: Reads GroupAssignment

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: GroupAssignment from StepBasic);
	---Purpose: Writes GroupAssignment

    Share (me; ent : GroupAssignment from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWGroupAssignment;
