-- File:	SWDRAW_ShapeTool.cdl
-- Created:	Tue Apr 22 18:34:27 1997
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


class ShapeTool  from SWDRAW 

    ---Purpose : Defines functions to control shapes (in way useful for XSTEP),
    --           additional features which should be basic, or call tools which
    --           are bound with transfer needs.           
    --           But these functions work on shapes, geometry, nothing else
    --           (no file, no model, no entity)


uses CString, Interpretor from Draw


is

    InitCommands (myclass; theCommands : in out Interpretor from Draw);
    ---Purpose : Defines and loads all basic functions for SWDRAW on Shapes

end ShapeTool;
