
-- File:	StepAP214_ApprovalItem.cdl
-- Created:	Tue Mar  9 17:02:25 1999
-- Author:	data exchange team
--		<det@androx.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class ApprovalItem from StepAP214 inherits SelectType from StepData


uses

    	AssemblyComponentUsageSubstitute from StepRepr,
	DocumentFile from StepBasic,
    	MaterialDesignation from StepRepr,
    	MechanicalDesignGeometricPresentationRepresentation from StepVisual,
	PresentationArea from StepVisual,
	Product from StepBasic,
	ProductDefinition from StepBasic,
	ProductDefinitionFormation from StepBasic,
	ProductDefinitionRelationship from StepBasic,
	PropertyDefinition from StepRepr,
	ShapeRepresentation from StepShape,
	SecurityClassification from StepBasic

is

	Create returns ApprovalItem;
	---Purpose : Returns a ApprovalItem SelectType

	CaseNum (me; ent : Transient) returns Integer is virtual;
	---Purpose: Recognizes a ApprovalItem Kind Entity that is :
    	--        1 -> AssemblyComponentUsageSubstitute
	--        2 -> DocumentFile
    	--        3 -> MaterialDesignation
    	--        4 -> MechanicalDesignGeometricPresentationRepresentation
	--        5 -> PresentationArea
    	--        6 -> Product
	--        7 -> ProductDefinition
    	--        8 -> ProductDefinitionFormation
	--        9 -> ProductDefinitionRelationship
	--        10 -> PropertyDefinition
    	--        11 -> ShapeRepresentation
	--        12 -> SecurityClassification
	--        0 else

    	AssemblyComponentUsageSubstitute (me) returns any AssemblyComponentUsageSubstitute is virtual ;
    	---Purpose : returns Value as a AssemblyComponentUsageSubstitute (Null if another type)
	
	DocumentFile (me) returns any DocumentFile is virtual;
	---Purpose : returns Value as a DocumentFile (Null if another type)
	
	MaterialDesignation (me) returns any MaterialDesignation is virtual;
	---Purpose : returns Value as a MaterialDesignation (Null if another type)
	
	MechanicalDesignGeometricPresentationRepresentation (me) returns any MechanicalDesignGeometricPresentationRepresentation is virtual;
	---Purpose : returns Value as a MechanicalDesignGeometricPresentationRepresentation (Null if another type)
	
	PresentationArea (me) returns any PresentationArea is virtual;
	---Purpose : returns Value as a PresentationArea (Null if another type)
	
	Product (me) returns any Product is virtual;
	---Purpose : returns Value as a Product (Null if another type)
	
	ProductDefinition (me) returns any ProductDefinition is virtual;
	---Purpose : returns Value as a ProductDefinition (Null if another type)
	
	ProductDefinitionFormation (me) returns any ProductDefinitionFormation is virtual;
	---Purpose : returns Value as a ProductDefinitionFormation (Null if another type)
	
	ProductDefinitionRelationship (me) returns any ProductDefinitionRelationship is virtual; 
	---Purpose : returns Value as aProductDefinitionRelationship (Null if another type)
	
	PropertyDefinition (me) returns any PropertyDefinition is virtual;
	---Purpose : returns Value as a PropertyDefinition (Null if another type)
	
	ShapeRepresentation (me) returns any ShapeRepresentation is virtual;
	---Purpose : returns Value as a ShapeRepresentation  (Null if another type)
	
	SecurityClassification (me) returns any SecurityClassification is virtual;
	---Purpose : returns Value as a SecurityClassification (Null if another type)
	
end ApprovalItem;
