-- File:	IntPoly_PntHasher.cdl
-- Created:	Tue Aug  8 11:32:21 1995
-- Author:	Stagiaire Alain JOURDAIN
--		<ajo@phobox>
---Copyright:	 Matra Datavision 1995


class PntHasher from IntPoly

uses  Pnt from gp

is    HashCode(myclass; Point : Pnt from gp;
                        Upper : Integer)
      returns Integer;
	---Purpose: Returns a HasCode value  for  the  Key <K>  in the
	--          range 0..Upper.
	---C++: inline
	
      IsEqual(myclass; Point1,Point2 : Pnt from gp)
      returns Boolean;
	---Purpose: Returns True  when the two  keys are the same. Two
	--          same  keys  must   have  the  same  hashcode,  the
	--          contrary is not necessary.
	---C++: inline
	
end PntHasher;
