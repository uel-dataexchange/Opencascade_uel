-- File:	RWStepVisual_RWExternallyDefinedCurveFont.cdl
-- Created:	Wed May 10 15:09:07 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWExternallyDefinedCurveFont from RWStepVisual

    ---Purpose: Read & Write tool for ExternallyDefinedCurveFont

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ExternallyDefinedCurveFont from StepVisual

is
    Create returns RWExternallyDefinedCurveFont from RWStepVisual;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ExternallyDefinedCurveFont from StepVisual);
	---Purpose: Reads ExternallyDefinedCurveFont

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ExternallyDefinedCurveFont from StepVisual);
	---Purpose: Writes ExternallyDefinedCurveFont

    Share (me; ent : ExternallyDefinedCurveFont from StepVisual;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWExternallyDefinedCurveFont;
