-- File:        AutoDesignDateAndTimeItem.cdl
-- Created:	Tue Mar  9 15:29:30 1999
-- Author:	data exchange team
--		<det@androx.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class PersonAndOrganizationItem from StepAP214 inherits ApprovalItem from StepAP214

	-- <PersonAndOrganizationItem> is an EXPRESS Select Type construct translation.
	-- it gathers : ApprovalPersonOrganization, AutoDesignDateAndPersonAssignment

uses

    	AppliedOrganizationAssignment from StepAP214
	
is

	Create returns PersonAndOrganizationItem;
	---Purpose : Returns a PersonAndOrganizationItem SelectType

	CaseNum (me; ent : Transient) returns Integer is redefined;
	---Purpose: Recognizes a APersonAndOrganizationItem Kind Entity that is :
    	--        1 -> AppliedOrganizationAssignment
    	--        2 -> AssemblyComponentUsageSubstitute
	--        3 -> DocumentFile
    	--        4 -> MaterialDesignation
    	--        5 -> MechanicalDesignGeometricPresentationRepresentation
	--        6 -> PresentationArea
    	--        7 -> Product
	--        8 -> ProductDefinition
    	--        9 -> ProductDefinitionFormation
	--    	  10 -> ProductDefinitionRelationship
	--        11 -> PropertyDefinition
    	--        12 -> ShapeRepresentation
    	--        13 -> SecurityClassification
	--        0 else


    	AppliedOrganizationAssignment (me) returns any AppliedOrganizationAssignment;
    	---Purpose : returns Value as a AppliedOrganizationAssignment (Null if another type)

	
end PersonAndOrganizationItem;
