-- File:	StepAP203_SpecifiedItem.cdl
-- Created:	Fri Nov 26 16:26:27 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class SpecifiedItem from StepAP203
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type SpecifiedItem

uses
    ProductDefinition from StepBasic,
    ShapeAspect from StepRepr

is
    Create returns SpecifiedItem from StepAP203;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of SpecifiedItem select type
	--          1 -> ProductDefinition from StepBasic
	--          2 -> ShapeAspect from StepRepr
	--          0 else

    ProductDefinition (me) returns ProductDefinition from StepBasic;
	---Purpose: Returns Value as ProductDefinition (or Null if another type)

    ShapeAspect (me) returns ShapeAspect from StepRepr;
	---Purpose: Returns Value as ShapeAspect (or Null if another type)

end SpecifiedItem;
