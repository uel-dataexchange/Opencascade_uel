-- File:	IGESDraw_ToolConnectPoint.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolConnectPoint  from IGESDraw

    ---Purpose : Tool to work on a ConnectPoint. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses ConnectPoint from IGESDraw,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolConnectPoint;
    ---Purpose : Returns a ToolConnectPoint, ready to work


    ReadOwnParams (me; ent : mutable ConnectPoint;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : ConnectPoint;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : ConnectPoint;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a ConnectPoint <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : ConnectPoint) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : ConnectPoint;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : ConnectPoint; entto : mutable ConnectPoint;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : ConnectPoint;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolConnectPoint;
