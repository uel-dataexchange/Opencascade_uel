-- File:        CsgShapeRepresentation.cdl
-- Created:     Mon Dec  4 12:02:25 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWCsgShapeRepresentation from RWStepShape

	---Purpose : Read & Write Module for CsgShapeRepresentation

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     CsgShapeRepresentation from StepShape,
     EntityIterator from Interface

is

	Create returns RWCsgShapeRepresentation;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable CsgShapeRepresentation from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : CsgShapeRepresentation from StepShape);

	Share(me; ent : CsgShapeRepresentation from StepShape; iter : in out EntityIterator);

end RWCsgShapeRepresentation;
