-- File:	BRepPrimAPI_MakeSphere.cdl
-- Created:	Thu Jul 22 19:23:53 1993
-- Author:	Remi LEQUETTE
--		<rle@nonox>
---Copyright:	 Matra Datavision 1993



class MakeSphere from BRepPrimAPI  inherits MakeOneAxis from BRepPrimAPI 

	---Purpose: Describes functions to build spheres or portions of spheres.
    	-- A MakeSphere object provides a framework for:
    	-- -   defining the construction of a sphere,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the result.

uses
    Pnt      from gp,
    Ax2      from gp,
    Sphere   from BRepPrim,
    OneAxis  from BRepPrim

raises
    DomainError from Standard

is
    Create(R : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public

    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(R, angle : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(R, angle1, angle2 : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(R, angle1, angle2, angle3 : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(Center : Pnt from gp; R : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(Center : Pnt from gp; R, angle : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(Center : Pnt from gp; R, angle1, angle2 : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(Center : Pnt from gp; R, angle1, angle2, angle3 : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(Axis : Ax2 from gp; R : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(Axis : Ax2 from gp; R, angle : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(Axis : Ax2 from gp; R, angle1, angle2 : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()

    Create(Axis : Ax2 from gp; R, angle1, angle2, angle3 : Real)
    returns MakeSphere from BRepPrimAPI
	---Purpose: Make a sphere of radius R.
	---Level: Public
    raises
    	DomainError from Standard; -- if R  <= Precision::Confusion()
    
    	---Purpose: For all algorithms The resulting shape is composed of
    	-- -   a lateral spherical face,
    	-- -   two planar faces parallel to the plane z = 0 if the
    	--   sphere is truncated in the v parametric direction, or
    	--   only one planar face if angle1 is equal to -p/2 or if
    	--     angle2 is equal to p/2 (these faces are circles in
    	--   case of a complete truncated sphere),
    	-- -   and in case of a portion of sphere, two planar faces
    	--   to shut the shape.(in the planes u = 0 and u = angle).   

    OneAxis(me : in out) returns Address;
	---Purpose: Returns the algorithm.
	---Level: Advanced

    Sphere(me : in out) returns Sphere from BRepPrim
	---Purpose: Returns the algorithm.
	--          
	---C++: return &
	---Level: Public 
    is static;

fields

    mySphere : Sphere from BRepPrim;

end MakeSphere;
