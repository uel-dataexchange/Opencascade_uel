-- File:        CurveStyleFontSelect.cdl
-- Created:     Fri Dec  1 11:11:11 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993



class CurveStyleFontSelect from StepVisual inherits SelectType from StepData

	-- <CurveStyleFontSelect> is an EXPRESS Select Type construct translation.
	-- it gathers : CurveStyleFont, PreDefinedCurveFont, ExternallyDefinedCurveFont

uses

	CurveStyleFont,
	PreDefinedCurveFont,
	ExternallyDefinedCurveFont
is

	Create returns CurveStyleFontSelect;
	---Purpose : Returns a CurveStyleFontSelect SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a CurveStyleFontSelect Kind Entity that is :
	--        1 -> CurveStyleFont
	--        2 -> PreDefinedCurveFont
	--        3 -> ExternallyDefinedCurveFont
	--        0 else

	CurveStyleFont (me) returns any CurveStyleFont;
	---Purpose : returns Value as a CurveStyleFont (Null if another type)

	PreDefinedCurveFont (me) returns any PreDefinedCurveFont;
	---Purpose : returns Value as a PreDefinedCurveFont (Null if another type)

	ExternallyDefinedCurveFont (me) returns any ExternallyDefinedCurveFont;
	---Purpose : returns Value as a ExternallyDefinedCurveFont (Null if another type)


end CurveStyleFontSelect;

