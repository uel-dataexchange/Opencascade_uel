-- File:	StepAP214_ExternallyDefinedClass.cdl
-- Created:	Wed May 10 15:09:06 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class ExternallyDefinedClass from StepAP214
inherits Class from StepAP214

    ---Purpose: Representation of STEP entity ExternallyDefinedClass

uses
    HAsciiString from TCollection,
    SourceItem from StepBasic,
    ExternalSource from StepBasic,
    ExternallyDefinedItem from StepBasic

is
    Create returns ExternallyDefinedClass from StepAP214;
	---Purpose: Empty constructor

    Init (me: mutable; aGroup_Name: HAsciiString from TCollection;
                       hasGroup_Description: Boolean;
                       aGroup_Description: HAsciiString from TCollection;
                       aExternallyDefinedItem_ItemId: SourceItem from StepBasic;
                       aExternallyDefinedItem_Source: ExternalSource from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    ExternallyDefinedItem (me) returns ExternallyDefinedItem from StepBasic;
	---Purpose: Returns data for supertype ExternallyDefinedItem
    SetExternallyDefinedItem (me: mutable; ExternallyDefinedItem: ExternallyDefinedItem from StepBasic);
	---Purpose: Set data for supertype ExternallyDefinedItem

fields
    theExternallyDefinedItem: ExternallyDefinedItem from StepBasic; -- supertype

end ExternallyDefinedClass;
