-- File:        OverRidingStyledItem.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWOverRidingStyledItem from RWStepVisual

	---Purpose : Read & Write Module for OverRidingStyledItem

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     OverRidingStyledItem from StepVisual,
     EntityIterator from Interface

is

	Create returns RWOverRidingStyledItem;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable OverRidingStyledItem from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : OverRidingStyledItem from StepVisual);

	Share(me; ent : OverRidingStyledItem from StepVisual; iter : in out EntityIterator);

end RWOverRidingStyledItem;
