-- File:	IGESDraw_ToolPlanar.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolPlanar  from IGESDraw

    ---Purpose : Tool to work on a Planar. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses Planar from IGESDraw,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolPlanar;
    ---Purpose : Returns a ToolPlanar, ready to work


    ReadOwnParams (me; ent : mutable Planar;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : Planar;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : Planar;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a Planar <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable Planar) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a Planar
    --           (NbMatrices forced to 1)

    DirChecker (me; ent : Planar) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : Planar;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : Planar; entto : mutable Planar;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : Planar;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolPlanar;
