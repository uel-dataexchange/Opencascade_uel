-- File:	StepGeom_GeomRepContextAndGlobUnitAssCtxAndGlobUncertaintyAssCtx.cdl
-- Created:	Thu Dec  7 14:45:21 1995
-- Author:	Frederic MAUPAS
--		<fma@pronox>
---Copyright:	 Matra Datavision 1995

class GeomRepContextAndGlobUnitAssCtxAndGlobUncertaintyAssCtx from StepGeom 

    inherits RepresentationContext from StepRepr

    -- This is a hand made implementation of EXPRESS ANDOR construct
    -- It gather 3 Types :
    -- 	      GeometricRepresentationContext
    -- 	      GlobalUnitAssignedContext
    -- 	      GlobalUncertaintyAssignedContext
    -- Common Supertype is RepresentationContext

uses 

    GeometricRepresentationContext      from StepGeom,
    GlobalUnitAssignedContext           from StepRepr,
    GlobalUncertaintyAssignedContext    from StepRepr,
    HArray1OfUncertaintyMeasureWithUnit from StepBasic,
    UncertaintyMeasureWithUnit          from StepBasic,
    HArray1OfNamedUnit                  from StepBasic, 
    NamedUnit                           from StepBasic,
    HAsciiString                        from TCollection, 
    Integer                             from Standard 


is

    Create returns mutable GeomRepContextAndGlobUnitAssCtxAndGlobUncertaintyAssCtx;
    
    Init (me : mutable;
          aContextIdentifier : mutable HAsciiString from TCollection;
          aContextType : mutable HAsciiString from TCollection) is redefined;

    Init(me : mutable;
         aContextIdentifier            : mutable HAsciiString                     from TCollection;
	 aContextType                  : mutable HAsciiString                     from TCollection;
	 aGeometricRepresentationCtx   : mutable GeometricRepresentationContext   from StepGeom;
	 aGlobalUnitAssignedCtx        : mutable GlobalUnitAssignedContext        from StepRepr;
    	 aGlobalUncertaintyAssignedCtx : mutable GlobalUncertaintyAssignedContext from StepRepr)
    is virtual;

    Init(me : mutable;
	 aContextIdentifier        : mutable HAsciiString                        from TCollection;
	 aContextType              : mutable HAsciiString                        from TCollection;
	 aCoordinateSpaceDimension : Integer                                     from Standard;
	 aUnits                    : mutable HArray1OfNamedUnit                  from StepBasic;
	 anUncertainty             : mutable HArray1OfUncertaintyMeasureWithUnit from StepBasic) 
    is virtual;

    -- ====================================== --
    -- Specific Methods for Field Data Access --
    -- ====================================== --

    SetGeometricRepresentationContext
    	(me : mutable; 
    	 aGeometricRepresentationContext : mutable GeometricRepresentationContext);

    GeometricRepresentationContext (me) 
    returns mutable GeometricRepresentationContext;

    SetGlobalUnitAssignedContext
    	(me : mutable; 
    	 aGlobalUnitAssignedContext : mutable GlobalUnitAssignedContext);

    GlobalUnitAssignedContext (me) 
    returns mutable GlobalUnitAssignedContext;

    SetGlobalUncertaintyAssignedContext
    	(me : mutable;
    	 aGlobalUncertaintyAssignedCtx : GlobalUncertaintyAssignedContext from StepRepr);
	 
    GlobalUncertaintyAssignedContext(me)
    returns GlobalUncertaintyAssignedContext from StepRepr;
    
    -- ============================================================================= --
    -- Specific Methods for ANDOR Field Data Access : GeometricRepresentationContext --
    -- ============================================================================= --
    
    SetCoordinateSpaceDimension(me : mutable; aCoordinateSpaceDimension : Integer);
    CoordinateSpaceDimension (me) returns Integer;

    -- ====================================================================== --
    -- Specific Methods for ANDOR Field Data Access GlobalUnitAssignedContext --
    -- ====================================================================== --

    SetUnits(me : mutable; aUnits : mutable HArray1OfNamedUnit);
    Units (me) returns mutable HArray1OfNamedUnit;
    UnitsValue (me; num : Integer) returns mutable NamedUnit;
    NbUnits (me) returns Integer;
	
    -- ============================================================================= --
    -- Specific Methods for ANDOR Field Data Access GlobalUncertaintyAssignedContext --
    -- ============================================================================= --

    SetUncertainty(me : mutable; aUncertainty : mutable HArray1OfUncertaintyMeasureWithUnit);
    Uncertainty (me) returns mutable HArray1OfUncertaintyMeasureWithUnit;
    UncertaintyValue (me; num : Integer) returns mutable UncertaintyMeasureWithUnit;
    NbUncertainty (me) returns Integer;

fields

    geometricRepresentationContext   : GeometricRepresentationContext   from StepGeom;
    globalUnitAssignedContext        : GlobalUnitAssignedContext        from StepRepr;
    globalUncertaintyAssignedContext : GlobalUncertaintyAssignedContext from StepRepr;

end GeomRepContextAndGlobUnitAssCtxAndGlobUncertaintyAssCtx;
