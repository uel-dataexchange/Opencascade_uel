-- File:        Date.cdl
-- Created:     Fri Dec  1 11:11:17 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class Date from StepBasic 

inherits TShared from MMgt

uses

	Integer from Standard
is

	Create returns mutable Date;
	---Purpose: Returns a Date

	Init (me : mutable;
	      aYearComponent : Integer from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetYearComponent(me : mutable; aYearComponent : Integer);
	YearComponent (me) returns Integer;

fields

	yearComponent : Integer from Standard;

end Date;
