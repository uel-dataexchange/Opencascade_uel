-- File:	IGESBasic_ToolSingularSubfigure.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolSingularSubfigure  from IGESBasic

    ---Purpose : Tool to work on a SingularSubfigure. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses SingularSubfigure from IGESBasic,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolSingularSubfigure;
    ---Purpose : Returns a ToolSingularSubfigure, ready to work


    ReadOwnParams (me; ent : mutable SingularSubfigure;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : SingularSubfigure;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : SingularSubfigure;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a SingularSubfigure <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : SingularSubfigure) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : SingularSubfigure;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : SingularSubfigure; entto : mutable SingularSubfigure;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : SingularSubfigure;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolSingularSubfigure;
