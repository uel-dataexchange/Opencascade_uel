-- File:	Image_Convertor.cdl
-- Created:	Wed Jul 28 16:08:03 1993
-- Author:	Jean Louis FRENKEL
--		<jlf@sparc3>
---Copyright:	 Matra Datavision 1993
    
    
class Convertor from Image

	---Purpose: This class is used to convert :
	--		a PseudoColorImage to a ColorImage
	--		a ColorImage to a PseudoColorImage
	--		a PseudoColorImage to a PseudoColorImage with a 
	--			different ColorMap.
	--
	--	    To convert a PseudoColoImage to a ColorImage we use
	--	    the PseudoColoImage ColorMap to compute the Color of each 
	--	    Image Pixel ( Lookup operation ) , the resulting image 
	--	    look similar as the original image.
	--
	--	    To convert a ColorImage to a PseudoColorImage or 
	--          a PseudoColorImage to another PseudoColorImage we use 
	--	    Dithering.
	--
	--	    A dither operation is an inverse lookup operation.For
	--	    example if we want to dither a ColorImage to a 
	--	    PseudoColorImage, for each Pixel in the ColorImage we search
	--	    in the PseudoColorImage ColorMap the Entry with the nearest
	--	    Color, then we write the ColorMap Entry Index in to the
	--	    PseudoColorImage. The result is a PseudoColorImage that when
	--	    it is displayed using its own ColorMap it will look as much 
	--          like the original ColorImage as possible.
	--
	--	    This class provides 2 Dithering method.
	--
	--	    DM_NearestColor : this dithering method is the simplest
	--	    one ,it just finds the nearest entry in the ColorMap.
	--	    This algorithm provide no provision for eliminating unwanted
	--	    contours in the dithered image.This algorithm is much 
	--	    faster on ColorRamp and ColorCube than on Generic
	--	    ColorMap.Indeed on ColorRamp and ColorCube ColorMap the
	--	    ColorMap Entry Index can be computed by using the ColorMap
	--	    BasePixel and ColorDimension.
	--	    
	--	    DM_ErrorDiffusion: In this method the difference ( error )
	--	    between the original and the dithered image is distribued
	--	    to the oginal image pixels immediatly to the right of and
	--	    below the last pixel processed. The ErrorDiffusion method
	--	    uses a "floyd-steinberg" error-distribution kernel.This
	--	    algorithm is fairly time-consuming, but can greatly reduce
	--	    contouring in the dithered image.
	--
    
uses
    ColorMap	 	from Aspect,
    GenericColorMap	from Aspect,
    ColorCubeColorMap	from Aspect,
    ColorRampColorMap	from Aspect,
    PseudoColorImage 	from Image,
    ColorImage 		from Image,
    DitheringMethod	from Image
    
is

    Create returns Convertor from Image;
	---Level: Public
	---Purpose: Create a Convertor object with the default DitheringMethod
	--	( DM_NearestColor ).

    SetDitheringMethod( me : in out ; 
			aMethod : in DitheringMethod from Image );
	---Level: Public
	---Purpose: Set DitheringMethod.

    Convert (me : in ;aColorImage: ColorImage from Image;
    	     		        aColorMap  : ColorMap from Aspect) 
    	returns mutable PseudoColorImage from Image;
	---Level: Public
	---Purpose: Dither a ColorImage into a PseudoColorImage using the
	--		 ColorMap parameter.
    
    Convert (me : in ; aPseudoColorImage: PseudoColorImage from Image;
    	     			 aColorMap	 : ColorMap from Aspect) 
    	returns mutable PseudoColorImage from Image;
	---Level: Public
	---Purpose: Dither a PseudoColorImage into a PseudoColorImage using the
	--		 ColorMap parameter.
    
    Convert (me : in; aPseudoColorImage: PseudoColorImage from Image)
    	returns mutable ColorImage from Image;
	---Level: Public
	---Purpose: Lookup a PseudoColorImage into a ColorImage using the
	--		PseudoColorImage ColorMap.

    --  *******************  Private Method   ******************* 

    NearestDithering(me : in; 
				aColorImage: ColorImage from Image ;
				aColorMap  : ColorMap   from Aspect) 
    	returns mutable PseudoColorImage from Image is private ;

    NearestDithering(me : in; 
			aPseudoColorImage : PseudoColorImage from Image ;
    	     		aColorMap	  : ColorMap   from Aspect) 
    	returns mutable PseudoColorImage from Image is private ;

    ErrorDiffusionDithering(me : in; 
			aColorImage       : ColorImage from Image ;
			aColorMap	  : ColorMap   from Aspect) 
    	returns mutable PseudoColorImage from Image is private ;

    ErrorDiffusionDithering(me : in; 
			aPseudoColorImage : PseudoColorImage from Image ;
			aColorMap	  : ColorMap   from Aspect) 
    	returns mutable PseudoColorImage from Image is private ;

fields

    myDitheringMethod : DitheringMethod from Image ;

end Convertor;
