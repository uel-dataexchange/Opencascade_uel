-- File:	StepToTopoDS_TranslateEdge.cdl
-- Created:	Fri Dec 16 14:48:04 1994
-- Author:	Frederic MAUPAS
--		<fma@stylox>
---Copyright:	 Matra Datavision 1994

class TranslateEdge from StepToTopoDS
    inherits Root from StepToTopoDS
    
    ---Purpose:
    --         

uses

    Edge               from StepShape,
    Tool               from StepToTopoDS,
    TranslateEdgeError from StepToTopoDS,
    Shape              from TopoDS,
    Edge               from TopoDS,
    Vertex             from TopoDS,
    Curve              from Geom2d,
    Surface            from Geom,
    EdgeCurve          from StepShape,
    Curve              from StepGeom,
    Vertex             from StepShape,
    Pcurve             from StepGeom,
    NMTool             from StepToTopoDS

raises NotDone from StdFail

is

    Create returns TranslateEdge;
    
    Create (E      : Edge from StepShape;
            T      : in out Tool from StepToTopoDS;
            NMTool : in out NMTool from StepToTopoDS)
    	returns TranslateEdge;
	    
    Init (me     : in out;
          E      : Edge from StepShape;
          T      : in out Tool from StepToTopoDS;
          NMTool : in out NMTool from StepToTopoDS);

    MakeFromCurve3D (me : in out; C3D : Curve from StepGeom;
    	    	     EC     : EdgeCurve from StepShape;        -- for messages
		     Vend   : Vertex from StepShape;      -- case of null edge
		     preci  : Real; E : in out Edge from TopoDS;
		     V1, V2 : in out Vertex from TopoDS;
		     T      : in out Tool from StepToTopoDS);
    ---Purpose:  Warning! C3D is assumed to be a Curve 3D ...
    --    other cases to checked before calling this

    MakePCurve (me; PCU : Pcurve from StepGeom; ConvSurf : Surface from Geom)
    	returns Curve from Geom2d;
    --  Null if failed

    Value (me) returns Shape from TopoDS
    	raises NotDone
	is static;
	---C++: return const &

    Error (me) returns TranslateEdgeError from StepToTopoDS;
    
fields

    myError  : TranslateEdgeError from StepToTopoDS;
    
    myResult : Shape              from TopoDS;
    
end TranslateEdge;
