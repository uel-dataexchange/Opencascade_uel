-- File:        ApprovalRelationship.cdl
-- Created:     Fri Dec  1 11:11:13 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class ApprovalRelationship from StepBasic 

inherits TShared from MMgt

uses

	HAsciiString from TCollection, 
	Approval from StepBasic
is

	Create returns mutable ApprovalRelationship;
	---Purpose: Returns a ApprovalRelationship

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aDescription : mutable HAsciiString from TCollection;
	      aRelatingApproval : mutable Approval from StepBasic;
	      aRelatedApproval : mutable Approval from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetName(me : mutable; aName : mutable HAsciiString);
	Name (me) returns mutable HAsciiString;
	SetDescription(me : mutable; aDescription : mutable HAsciiString);
	Description (me) returns mutable HAsciiString;
	SetRelatingApproval(me : mutable; aRelatingApproval : mutable Approval);
	RelatingApproval (me) returns mutable Approval;
	SetRelatedApproval(me : mutable; aRelatedApproval : mutable Approval);
	RelatedApproval (me) returns mutable Approval;

fields

	name : HAsciiString from TCollection;
	description : HAsciiString from TCollection;
	relatingApproval : Approval from StepBasic;
	relatedApproval : Approval from StepBasic;

end ApprovalRelationship;
