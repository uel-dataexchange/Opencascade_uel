-- File:        CoordinatedUniversalTimeOffset.cdl
-- Created:     Fri Dec  1 11:11:17 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class CoordinatedUniversalTimeOffset from StepBasic 

inherits TShared from MMgt

uses

	Integer from Standard, 
	AheadOrBehind from StepBasic, 
	Boolean from Standard
is

	Create returns mutable CoordinatedUniversalTimeOffset;
	---Purpose: Returns a CoordinatedUniversalTimeOffset

	Init (me : mutable;
	      aHourOffset : Integer from Standard;
	      hasAminuteOffset : Boolean from Standard;
	      aMinuteOffset : Integer from Standard;
	      aSense : AheadOrBehind from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetHourOffset(me : mutable; aHourOffset : Integer);
	HourOffset (me) returns Integer;
	SetMinuteOffset(me : mutable; aMinuteOffset : Integer);
	UnSetMinuteOffset (me:mutable);
	MinuteOffset (me) returns Integer;
	HasMinuteOffset (me) returns Boolean;
	SetSense(me : mutable; aSense : AheadOrBehind);
	Sense (me) returns AheadOrBehind;

fields

	hourOffset : Integer from Standard;
	minuteOffset : Integer from Standard;   -- OPTIONAL can be NULL
	sense : AheadOrBehind from StepBasic; -- an Enumeration
	hasMinuteOffset : Boolean from Standard;

end CoordinatedUniversalTimeOffset;
