-- File:        BRepBlend_HCurveToolGen.cdl
-- Created:	Mon Jul 17 16:25:23 1995
-- Author:	Laurent BUCHARD
--		<lbr@mastox>
---Copyright:	 Matra Datavision 1995


generic class HCurveToolGen from BRepBlend (
     CurveGen  as any)

uses 
     Array1OfReal    from TColStd,
     Shape           from GeomAbs,
     CurveType       from GeomAbs,
     Vec             from gp,
     Pnt             from gp,
     Circ            from gp,
     Elips           from gp,
     Hypr            from gp,
     Parab           from gp,
     Lin             from gp,
     BezierCurve     from Geom,
     BSplineCurve    from Geom
     
raises
    
    OutOfRange          from Standard,
    NoSuchObject        from Standard,
    DomainError         from Standard
 
is

    --
    --     Global methods - Apply to the whole curve.
    --     
    
    FirstParameter(myclass; C: CurveGen) returns Real
    	---C++: inline
    ;
    

    LastParameter(myclass; C: CurveGen) returns Real
    	---C++: inline    
    ;

    --
    -- Services to break the curves to the expected continuity
    -- 
    --  If  for example you  need the  curve to  be C2  and the method
    --  Continuity   returns you something lower than   C2 (say C1 for
    --  example).
    --  
    --  First  compute the   number  of intervals  with  the requested
    --  continuity with the method  NbIntervals().   Note that if  the
    --  continuity  is higher than the one   you need NbIntervals will
    --  return 1.
    --  
    --  Then you get the parameters  bounding  the intervals with  the
    --  method  Intervals,   using   an array    of  length  at  least
    --  NbIntervals()+1.
    -- 
    -- If you need  to create a curve  with a restricted span you  can
    -- use the method Trim().

    
    Continuity(myclass; C: CurveGen) returns Shape from GeomAbs
	---Purpose: 
	---C++: inline
    ;
    
    NbIntervals(myclass; C: CurveGen; S : Shape from GeomAbs) returns Integer
	---Purpose: Returns  the number  of  intervals for  continuity
	--          <S>. May be one if Continuity(myclass) >= <S>
	---C++: inline
    ;
    
    Intervals(myclass; C: CurveGen; T : in out Array1OfReal from TColStd; 
    	          S : Shape from GeomAbs)
	---Purpose: Stores in <T> the  parameters bounding the intervals
	--          of continuity <S>.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
    raises
    	OutOfRange from Standard
    ---C++: inline
    ;
    
    IsClosed(myclass; C: CurveGen) returns Boolean
    ---C++: inline    
    ;
     
    IsPeriodic(myclass; C: CurveGen) returns Boolean
    ---C++: inline
    ;
    
    Period(myclass; C: CurveGen) returns Real
    raises
    	DomainError from Standard -- if the curve is not periodic
    ---C++: inline	
    ;
     
    Value(myclass; C: CurveGen; U : Real) returns Pnt from gp
         --- Purpose : Computes the point of parameter U on the curve.
    ---C++: inline
    ;
    
    D0 (myclass; C: CurveGen; U : Real; P : out Pnt from gp)
         --- Purpose : Computes the point of parameter U on the curve.
    ---C++: inline
    ;
    
    D1 (myclass; C: CurveGen; U : Real; P : out Pnt from gp ; V : out Vec from gp)
         --- Purpose : Computes the point of parameter U on the curve with its
         --  first derivative.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C1.
    ---C++: inline
    ;
    
    D2 (myclass; C: CurveGen; U : Real; P : out Pnt from gp; V1, V2 : out Vec from gp)
        --- Purpose :
        --  Returns the point P of parameter U, the first and second
        --  derivatives V1 and V2.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C2.
    ---C++: inline
     ;

    D3 (myclass; C: CurveGen; U : Real; P : out Pnt from gp; V1, V2, V3 : out Vec from gp)
        --- Purpose :
        --  Returns the point P of parameter U, the first, the second 
        --  and the third derivative.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C3.
    ---C++: inline
     ;
        
    DN (myclass; C: CurveGen; U : Real; N : Integer)   returns Vec from gp
        --- Purpose :
        --  The returned vector gives the value of the derivative for the 
        --  order of derivation N.
     raises  
    	DomainError from Standard,
        --- Purpose : Raised if the continuity of the current interval
        --  is not CN.
        OutOfRange from Standard
        --- Purpose : Raised if N < 1.            
    ---C++: inline
     ;

    Resolution(myclass; C: CurveGen; R3d : Real) returns Real
         ---Purpose :  Returns the parametric  resolution corresponding
         --         to the real space resolution <R3d>.
    ---C++: inline
    ;   
        
    GetType(myclass; C: CurveGen) returns CurveType from GeomAbs
	---Purpose: Returns  the  type of the   curve  in the  current
	--          interval :   Line,   Circle,   Ellipse, Hyperbola,
	--          Parabola, BezierCurve, BSplineCurve, OtherCurve.
    ---C++: inline
    ;

    --
    --     The following methods must  be called when GetType returned
    --     the corresponding type.
    --     

     Line(myclass; C: CurveGen) returns Lin from gp
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;
     
     Circle(myclass; C: CurveGen) returns Circ from gp
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;
     
     Ellipse(myclass; C: CurveGen) returns Elips from gp
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;
     
     Hyperbola(myclass; C: CurveGen) returns  Hypr from gp
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;
     
     Parabola(myclass; C: CurveGen) returns Parab from gp
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;
     
     Bezier(myclass; C: CurveGen) returns BezierCurve from Geom
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;
    
     BSpline(myclass; C: CurveGen) returns BSplineCurve from Geom
     raises 
    	NoSuchObject from Standard
    ---C++: inline
     ;

    



    NbSamples(myclass; C: CurveGen; U0,U1: Real from Standard) 
    returns Integer from Standard;

end HCurveToolGen;


