-- File:	AppCont_Function.cdl
-- Created:	Wed Sep  1 15:17:55 1993
-- Author:	Laurent PAINNOT
--		<lpa@nonox>
---Copyright:	 Matra Datavision 1993


deferred class Function from AppCont

    ---Purpose: deferred class describing a continous 3d function f(u)


uses Pnt from gp,
     Vec from gp

is

    Delete(me:out) is virtual;
    ---C++: alias "Standard_EXPORT virtual ~AppCont_Function(){Delete() ; }"
    

    FirstParameter(me) returns Real
    	---Purpose: returns the first parameter of the function.
    is deferred;

    LastParameter(me) returns Real
    	---Purpose: returns the last parameter of the function.
    is deferred;

    Value(me; U: Real) returns Pnt
    	---Purpose: returns the point at parameter <U>.
    is deferred;

    D1(me; U: Real; P: in out Pnt; V: in out Vec) returns Boolean
    	---Purpose: returns the point and the derivative values at
    	--          the parameter <U>.
    is deferred;
    
    
end Function;    
