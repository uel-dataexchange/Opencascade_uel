-- File:	RWStepBasic_RWVersionedActionRequest.cdl
-- Created:	Fri Nov 26 16:26:40 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWVersionedActionRequest from RWStepBasic

    ---Purpose: Read & Write tool for VersionedActionRequest

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    VersionedActionRequest from StepBasic

is
    Create returns RWVersionedActionRequest from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : VersionedActionRequest from StepBasic);
	---Purpose: Reads VersionedActionRequest

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: VersionedActionRequest from StepBasic);
	---Purpose: Writes VersionedActionRequest

    Share (me; ent : VersionedActionRequest from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWVersionedActionRequest;
