-- File:        ConversionBasedUnitAndPlaneAngleUnit.cdl
-- Created:     Mon Dec  4 12:02:37 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWConversionBasedUnitAndPlaneAngleUnit from RWStepBasic

	---Purpose : Read & Write Module for ConversionBasedUnitAndPlaneAngleUnit

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ConversionBasedUnitAndPlaneAngleUnit from StepBasic,
     EntityIterator from Interface

is

	Create returns RWConversionBasedUnitAndPlaneAngleUnit;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ConversionBasedUnitAndPlaneAngleUnit from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : ConversionBasedUnitAndPlaneAngleUnit from StepBasic);

	Share(me; ent : ConversionBasedUnitAndPlaneAngleUnit from StepBasic; iter : in out EntityIterator);

end RWConversionBasedUnitAndPlaneAngleUnit;
