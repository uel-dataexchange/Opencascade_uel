-- File:        PresentationLayerAssignment.cdl
-- Created:     Mon Dec  4 12:02:29 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPresentationLayerAssignment from RWStepVisual

	---Purpose : Read & Write Module for PresentationLayerAssignment

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PresentationLayerAssignment from StepVisual,
     EntityIterator from Interface

is

	Create returns RWPresentationLayerAssignment;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PresentationLayerAssignment from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : PresentationLayerAssignment from StepVisual);

	Share(me; ent : PresentationLayerAssignment from StepVisual; iter : in out EntityIterator);

end RWPresentationLayerAssignment;
