-- File:	StepAP203_PersonOrganizationItem.cdl
-- Created:	Fri Nov 26 16:26:27 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class PersonOrganizationItem from StepAP203
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type PersonOrganizationItem

uses
    Change from StepAP203,
    StartWork from StepAP203,
    ChangeRequest from StepAP203,
    StartRequest from StepAP203,
    ConfigurationItem from StepRepr,
    Product from StepBasic,
    ProductDefinitionFormation from StepBasic,
    ProductDefinition from StepBasic,
    Contract from StepBasic,
    SecurityClassification from StepBasic

is
    Create returns PersonOrganizationItem from StepAP203;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of PersonOrganizationItem select type
	--          1 -> Change from StepAP203
	--          2 -> StartWork from StepAP203
	--          3 -> ChangeRequest from StepAP203
	--          4 -> StartRequest from StepAP203
	--          5 -> ConfigurationItem from StepRepr
	--          6 -> Product from StepBasic
	--          7 -> ProductDefinitionFormation from StepBasic
	--          8 -> ProductDefinition from StepBasic
	--          9 -> Contract from StepBasic
	--          10 -> SecurityClassification from StepBasic
	--          0 else

    Change (me) returns Change from StepAP203;
	---Purpose: Returns Value as Change (or Null if another type)

    StartWork (me) returns StartWork from StepAP203;
	---Purpose: Returns Value as StartWork (or Null if another type)

    ChangeRequest (me) returns ChangeRequest from StepAP203;
	---Purpose: Returns Value as ChangeRequest (or Null if another type)

    StartRequest (me) returns StartRequest from StepAP203;
	---Purpose: Returns Value as StartRequest (or Null if another type)

    ConfigurationItem (me) returns ConfigurationItem from StepRepr;
	---Purpose: Returns Value as ConfigurationItem (or Null if another type)

    Product (me) returns Product from StepBasic;
	---Purpose: Returns Value as Product (or Null if another type)

    ProductDefinitionFormation (me) returns ProductDefinitionFormation from StepBasic;
	---Purpose: Returns Value as ProductDefinitionFormation (or Null if another type)

    ProductDefinition (me) returns ProductDefinition from StepBasic;
	---Purpose: Returns Value as ProductDefinition (or Null if another type)

    Contract (me) returns Contract from StepBasic;
	---Purpose: Returns Value as Contract (or Null if another type)

    SecurityClassification (me) returns SecurityClassification from StepBasic;
	---Purpose: Returns Value as SecurityClassification (or Null if another type)

end PersonOrganizationItem;
