-- File:	RWStepDimTol_RWDatumReference.cdl
-- Created:	Wed Jun  4 13:34:35 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWDatumReference from RWStepDimTol

    ---Purpose: Read & Write tool for DatumReference

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    DatumReference from StepDimTol

is
    Create returns RWDatumReference from RWStepDimTol;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : DatumReference from StepDimTol);
	---Purpose: Reads DatumReference

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: DatumReference from StepDimTol);
	---Purpose: Writes DatumReference

    Share (me; ent : DatumReference from StepDimTol;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWDatumReference;
