-- File:	StepGeom_OrientedSurface.cdl
-- Created:	Fri Jan  4 17:42:44 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class OrientedSurface from StepGeom
inherits Surface from StepGeom

    ---Purpose: Representation of STEP entity OrientedSurface

uses
    HAsciiString from TCollection

is
    Create returns OrientedSurface from StepGeom;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aOrientation: Boolean);
	---Purpose: Initialize all fields (own and inherited)

    Orientation (me) returns Boolean;
	---Purpose: Returns field Orientation
    SetOrientation (me: mutable; Orientation: Boolean);
	---Purpose: Set field Orientation

fields
    theOrientation: Boolean;

end OrientedSurface;
