-- File:        ApplicationProtocolDefinition.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWApplicationProtocolDefinition from RWStepBasic

	---Purpose : Read & Write Module for ApplicationProtocolDefinition

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ApplicationProtocolDefinition from StepBasic,
     EntityIterator from Interface

is

	Create returns RWApplicationProtocolDefinition;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ApplicationProtocolDefinition from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : ApplicationProtocolDefinition from StepBasic);

	Share(me; ent : ApplicationProtocolDefinition from StepBasic; iter : in out EntityIterator);

end RWApplicationProtocolDefinition;
