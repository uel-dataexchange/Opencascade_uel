-- File:        DateAndTime.cdl
-- Created:     Mon Dec  4 12:02:25 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWDateAndTime from RWStepBasic

	---Purpose : Read & Write Module for DateAndTime

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     DateAndTime from StepBasic,
     EntityIterator from Interface

is

	Create returns RWDateAndTime;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable DateAndTime from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : DateAndTime from StepBasic);

	Share(me; ent : DateAndTime from StepBasic; iter : in out EntityIterator);

end RWDateAndTime;
