-- File:	IGESSolid_ToolSphere.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolSphere  from IGESSolid

    ---Purpose : Tool to work on a Sphere. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses Sphere from IGESSolid,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolSphere;
    ---Purpose : Returns a ToolSphere, ready to work


    ReadOwnParams (me; ent : mutable Sphere;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : Sphere;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : Sphere;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a Sphere <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : Sphere) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : Sphere;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : Sphere; entto : mutable Sphere;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : Sphere;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolSphere;
