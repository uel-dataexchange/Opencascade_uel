-- File:	StepData_SelectInt.cdl
-- Created:	Mon Dec 16 16:23:07 1996
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996


class SelectInt  from StepData    inherits SelectMember

    ---Purpose : A SelectInt is a SelectMember specialised for a basic integer
    --           type in a select which also accepts entities : this one has
    --           NO NAME.
    --           For a named select, see SelectNamed

uses CString, Logical

is

    Create returns mutable SelectInt;

    Kind (me) returns Integer  is redefined;
    --  possible kind for Int : integer boolean logical enum(without text)

    SetKind  (me : mutable; kind : Integer)  is redefined;
    --  called by various Set*

    Int  (me) returns Integer  is redefined;

    SetInt (me : mutable; val : Integer)  is redefined;

fields

    thekind : Integer;
    theval  : Integer;

end SelectInt;
