-- File:	Storage_Root.cdl
-- Created:	Mon Feb 24 16:30:08 1997
-- Author:	Kernel
--		<kernel@parigox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997

class Root from Storage

inherits TShared from MMgt 
    	---Purpose:
    	-- A root object extracted from a Storage_Data object.
    	-- A Storage_Root encapsulates a persistent
    	-- object which is a root of a Storage_Data object.
    	-- It contains additional information: the name and
    	-- the data type of the persistent object.
    	-- When retrieving a Storage_Data object from a
    	-- container (for example, a file) you access its
    	-- roots with the function Roots which returns a
    	-- sequence of root objects. The provided functions
    	-- allow you to request information about each root of the sequence.
    	-- You do not create explicit roots: when inserting
    	-- data in a Storage_Data object, you just provide
    	-- the persistent object and optionally its name to the function AddRoot.
uses AsciiString from TCollection

is
    Create returns mutable Root from Storage;

    Create(aName    : AsciiString from TCollection;
    	   anObject : Persistent  from Standard) returns mutable Root from Storage;

    SetName(me : mutable; aName    : AsciiString from TCollection);
    Name(me) returns AsciiString from TCollection;
    	---Purpose:
    	-- Returns the name of this root object.
    	--   The name may have been given explicitly when
    	-- the root was inserted into the Storage_Data
    	-- object. If not, the name is a reference number
    	-- which was assigned automatically by the driver
    	-- when writing the set of data into the container.
    	-- When naming the roots, it is easier to retrieve
    	-- objects by significant references rather than by
    	-- references without any semantic values.
    	-- Warning
    	-- The returned string will be empty if you call this
    	-- function before having named this root object,
    	-- either explicitly, or when writing the set of data
    	-- into the container.    
    
    SetObject(me : mutable; anObject : Persistent  from Standard);
    Object(me) returns mutable Persistent  from Standard;
    	---Purpose:
    	-- Returns the persistent object encapsulated by this root.    
    Type(me) returns AsciiString from TCollection;
    	---Purpose: Returns the name of this root type.   
    
    SetReference(me : mutable; aRef : Integer from Standard) is private;
    Reference(me) returns Integer from Standard is private;
    SetType(me : mutable; aType : AsciiString from TCollection) is private;
    
    fields
    	
    	myName   : AsciiString from TCollection;
	myType   : AsciiString from TCollection;
	myObject : Persistent  from Standard;
	myRef    : Integer     from Standard;
	
    friends class Schema from Storage
    
end;
