-- File:        BezierSurface.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWBezierSurface from RWStepGeom

	---Purpose : Read & Write Module for BezierSurface

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     BezierSurface from StepGeom,
     EntityIterator from Interface

is

	Create returns RWBezierSurface;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable BezierSurface from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : BezierSurface from StepGeom);

	Share(me; ent : BezierSurface from StepGeom; iter : in out EntityIterator);

end RWBezierSurface;
