-- File:	StepFEA_DegreeOfFreedom.cdl
-- Created:	Sat Dec 14 11:02:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class DegreeOfFreedom from StepFEA
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type DegreeOfFreedom

uses
    SelectMember from StepData,
    EnumeratedDegreeOfFreedom from StepFEA,
    HAsciiString from TCollection

is
    Create returns DegreeOfFreedom from StepFEA;
	---Purpose: Empty constructor
	
    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of CurveElementFreedom select type
	--          return 0

    CaseMem (me; ent: SelectMember from StepData) returns Integer is redefined;
	---Purpose: Recognizes a items of select member CurveElementFreedomMember
	--          1 -> EnumeratedCurveElementFreedom
	--          2 -> ApplicationDefinedDegreeOfFreedom
	--          0 else
	
    NewMember(me) returns SelectMember from StepData is redefined;
	---Purpose: Returns a new select member the type CurveElementFreedomMember

    SetEnumeratedDegreeOfFreedom (me:in out; aVal: EnumeratedDegreeOfFreedom from StepFEA);
	---Purpose: Returns Value as EnumeratedDegreeOfFreedom (or Null if another type)
	
    EnumeratedDegreeOfFreedom (me) returns EnumeratedDegreeOfFreedom from StepFEA;
    	---Purpose: Returns Value as EnumeratedDegreeOfFreedom (or Null if another type)
	
    SetApplicationDefinedDegreeOfFreedom(me: in out; aVal :HAsciiString from TCollection);
	---Purpose: Set Value for ApplicationDefinedDegreeOfFreedom

    ApplicationDefinedDegreeOfFreedom (me) returns HAsciiString from TCollection;
	---Purpose: Returns Value as ApplicationDefinedDegreeOfFreedom (or Null if another type)

end DegreeOfFreedom;
