-- File:	Graphic3d_Texture1Dsegment.cdl
-- Created:	Mon Jul 28 10:40:23 1997
-- Author:	Pierre CHALAMET
--		<pct@sgi93>
---Copyright:	 Matra Datavision 1997 

class  Texture1Dsegment  from  Graphic3d 
    
inherits  Texture1D  from  Graphic3d  

 
    ---Purpose:  This class provides the implementation
    -- of a 1D texture applyable along a segment.
    -- You might use the SetSegment() method
    -- to set the way the texture is "streched" on facets. 


uses 
    NameOfTexture1D  from  Graphic3d, 
    StructureManager      from  Graphic3d 

is 
    Create(VM  :  StructureManager  from  Graphic3d; 
    	   FileName  :  CString  from  Standard)  returns  mutable  Texture1Dsegment  from  Graphic3d; 
    ---Purpose: Creates a texture from a file


    Create(VM  :  StructureManager  from  Graphic3d; 
    	   NOT  :  NameOfTexture1D  from  Graphic3d)  returns  mutable  Texture1Dsegment  from  Graphic3d;  
    ---Purpose: Creates a texture from a predefined texture name set.
     
    SetSegment(me  :  mutable; 
    	       X1,Y1,Z1  :  ShortReal  from  Standard; 
	       X2,Y2,Z2  :  ShortReal  from  Standard);
    ---Purpose: Sets the texture application bounds. Defines the way
    -- the texture is stretched across facets.
    -- Default values are <0.0, 0.0, 0.0> , <0.0, 0.0, 1.0>

  
    --
    -- inquire methods
    --
    Segment(me;
            X1,Y1,Z1, X2,Y2,Z2 : out ShortReal from Standard);
    ---Purpose: Returns the values of the current segment X1, Y1, Z1 , X2, Y2, Z2.
    
fields    
    MyX1,MyY1,MyZ1  :  ShortReal  from  Standard; 
    MyX2,MyY2,MyZ2  :  ShortReal  from  Standard;
      
end  Texture1Dsegment; 

