-- File:	StepBasic_Document.cdl
-- Created:	Thu May 11 16:38:00 2000 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class Document from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity Document

uses
    HAsciiString from TCollection,
    DocumentType from StepBasic

is
    Create returns Document from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aId: HAsciiString from TCollection;
                       aName: HAsciiString from TCollection;
                       hasDescription: Boolean;
                       aDescription: HAsciiString from TCollection;
                       aKind: DocumentType from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Id (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Id
    SetId (me: mutable; Id: HAsciiString from TCollection);
	---Purpose: Set field Id

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description
    HasDescription (me) returns Boolean;
	---Purpose: Returns True if optional field Description is defined

    Kind (me) returns DocumentType from StepBasic;
	---Purpose: Returns field Kind
    SetKind (me: mutable; Kind: DocumentType from StepBasic);
	---Purpose: Set field Kind

fields
    theId: HAsciiString from TCollection;
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection; -- optional
    theKind: DocumentType from StepBasic;
    defDescription: Boolean; -- flag "is Description defined"

end Document;
