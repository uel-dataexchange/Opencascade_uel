-- File:	BOP_SolidSolidHistoryCollector.cdl
-- Created:	Thu Mar 20 15:39:35 2003
-- Author:	Michael KLOKOV
--		<mkk@kurox>
---Copyright:	Open CASCADE 2003

class SolidSolidHistoryCollector from BOP 
    inherits HistoryCollector from BOP

uses
    Shape from TopoDS,
    Operation from BOP,
    PDSFiller from BOPTools,
    ListOfShape from TopTools
is
    Create(theShape1   : Shape from TopoDS;
    	   theShape2   : Shape from TopoDS;
	   theOperation: Operation from BOP)
    	returns SolidSolidHistoryCollector from BOP;

    AddNewShape(me: mutable; theOldShape: Shape from TopoDS;
    	    	    	    theNewShape: Shape from TopoDS;
    	    	    	    theDSFiller: PDSFiller from BOPTools);

    SetResult(me: mutable; theResult: Shape from TopoDS;
    	    	    	   theDSFiller: PDSFiller from BOPTools)
    	is redefined virtual;

end SolidSolidHistoryCollector from BOP;
