-- File:	RWStepDimTol_RWTotalRunoutTolerance.cdl
-- Created:	Wed Jun  4 13:34:34 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWTotalRunoutTolerance from RWStepDimTol

    ---Purpose: Read & Write tool for TotalRunoutTolerance

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    TotalRunoutTolerance from StepDimTol

is
    Create returns RWTotalRunoutTolerance from RWStepDimTol;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : TotalRunoutTolerance from StepDimTol);
	---Purpose: Reads TotalRunoutTolerance

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: TotalRunoutTolerance from StepDimTol);
	---Purpose: Writes TotalRunoutTolerance

    Share (me; ent : TotalRunoutTolerance from StepDimTol;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWTotalRunoutTolerance;
