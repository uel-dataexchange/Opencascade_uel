-- File:	XSControl_SelectForTransfer.cdl
-- Created:	Tue Mar 26 14:03:27 1996
-- Author:	Christian CAILLET
--		<cky@fidox>
---Copyright:	 Matra Datavision 1996


class SelectForTransfer  from XSControl   inherits SelectExtract  from IFSelect

    ---Purpose : This selection selects the entities which are recognised for
    --           transfer by an Actor for Read : current one or another one.
    --           
    --           An Actor is an operator which runs transfers from interface
    --           entities to objects for Imagine. It has a method to recognize
    --           the entities it can process (by default, it recognises all,
    --           this method can be redefined).
    --           
    --           A TransferReader brings an Actor, according to the currently
    --           selected norm and transfer conditions.
    --           
    --           This selection considers, either the current Actor (brought by
    --           the TransferReader, updated as required), or a precise one.

uses AsciiString from TCollection, InterfaceModel,
     ActorOfTransientProcess, TransferReader

is

    Create returns mutable SelectForTransfer;
    ---Purpose : Creates a SelectForTransfer, non initialised
    --           it sorts nothing, unless an Actor has been defined

    Create (TR : TransferReader) returns mutable SelectForTransfer;
    ---Purpose : Creates a SelectForTransfer, which will work with the
    --           currently defined Actor brought by the TransferReader

    SetReader (me : mutable; TR : TransferReader);
    ---Purpose : Sets a TransferReader to sort entities : it brings the Actor,
    --           which may change, while the TransferReader does not

    SetActor (me : mutable; act : mutable ActorOfTransientProcess);
    ---Purpose : Sets a precise actor to sort entities
    --           This definition oversedes the creation with a TransferReader

    Actor (me) returns ActorOfTransientProcess;
    ---Purpose : Returns the Actor used as precised one.
    --           Returns a Null Handle for a creation from a TransferReader
    --           without any further setting

    Reader (me) returns TransferReader;
    ---Purpose : Returns the Reader (if created with a Reader)
    --           Returns a Null Handle if not created with a Reader


    Sort (me; rank : Integer; ent : Transient; model : InterfaceModel)
        returns Boolean;
    ---Purpose : Returns True for an Entity which is recognized by the Actor,
    --           either the precised one, or the one defined by TransferReader
     
    --Sort (me;  ent : in out Transient) returns Boolean;
     
    ExtractLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium : "Recognized for Transfer [(current actor)]"

fields

    theTR : TransferReader;
    theAC : ActorOfTransientProcess;

end SelectForTransfer;
