-- File:	IGESSolid_ToolEdgeList.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolEdgeList  from IGESSolid

    ---Purpose : Tool to work on a EdgeList. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses EdgeList from IGESSolid,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolEdgeList;
    ---Purpose : Returns a ToolEdgeList, ready to work


    ReadOwnParams (me; ent : mutable EdgeList;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : EdgeList;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : EdgeList;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a EdgeList <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : EdgeList) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : EdgeList;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : EdgeList; entto : mutable EdgeList;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : EdgeList;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolEdgeList;
