-- File:        ShapeAspect.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWShapeAspect from RWStepRepr

	---Purpose : Read & Write Module for ShapeAspect

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ShapeAspect from StepRepr,
     EntityIterator from Interface

is

	Create returns RWShapeAspect;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ShapeAspect from StepRepr);

	WriteStep (me; SW : in out StepWriter; ent : ShapeAspect from StepRepr);

	Share(me; ent : ShapeAspect from StepRepr; iter : in out EntityIterator);

end RWShapeAspect;
