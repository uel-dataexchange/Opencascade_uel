-- File:        Face.cdl
-- Created:     Fri Dec  1 11:11:20 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class Face from StepShape 

inherits TopologicalRepresentationItem from StepShape 

uses

	HArray1OfFaceBound from StepShape, 
	FaceBound from StepShape, 
	HAsciiString from TCollection
is

	Create returns mutable Face;
	---Purpose: Returns a Face


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aBounds : mutable HArray1OfFaceBound from StepShape) is virtual;

	-- Specific Methods for Field Data Access --

	SetBounds(me : mutable; aBounds : mutable HArray1OfFaceBound)
    	is virtual;
	Bounds (me) returns mutable HArray1OfFaceBound
    	is virtual;
	BoundsValue (me; num : Integer) returns mutable FaceBound
    	is virtual;
	NbBounds (me) returns Integer
    	is virtual;

fields

	bounds : HArray1OfFaceBound from StepShape;

end Face;
