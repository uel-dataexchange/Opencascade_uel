-- File:        StyledItem.cdl
-- Created:     Fri Dec  1 11:11:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class StyledItem from StepVisual 

inherits RepresentationItem from StepRepr

uses

	HArray1OfPresentationStyleAssignment from StepVisual, 
	PresentationStyleAssignment from StepVisual, 
	HAsciiString from TCollection
is

	Create returns mutable StyledItem;
	---Purpose: Returns a StyledItem


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aStyles : mutable HArray1OfPresentationStyleAssignment from StepVisual;
	      aItem : mutable RepresentationItem from StepRepr) is virtual;

	-- Specific Methods for Field Data Access --

	SetStyles(me : mutable; aStyles : mutable HArray1OfPresentationStyleAssignment);
	Styles (me) returns mutable HArray1OfPresentationStyleAssignment;
	StylesValue (me; num : Integer) returns mutable PresentationStyleAssignment;
	NbStyles (me) returns Integer;
	SetItem(me : mutable; aItem : mutable RepresentationItem);
	Item (me) returns mutable RepresentationItem;

fields

	styles : HArray1OfPresentationStyleAssignment from StepVisual;
	item : RepresentationItem from StepRepr;

end StyledItem;
