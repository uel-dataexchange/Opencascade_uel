-- File:        SolidAngleMeasureWithUnit.cdl
-- Created:     Fri Dec  1 11:11:27 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class SolidAngleMeasureWithUnit from StepBasic 

inherits MeasureWithUnit from StepBasic 

uses

	Real from Standard, 
	NamedUnit from StepBasic
is

	Create returns mutable SolidAngleMeasureWithUnit;
	---Purpose: Returns a SolidAngleMeasureWithUnit


end SolidAngleMeasureWithUnit;
