-- File:	RWStepFEA_RWFeaSecantCoefficientOfLinearThermalExpansion.cdl
-- Created:	Thu Dec 12 17:51:06 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFeaSecantCoefficientOfLinearThermalExpansion from RWStepFEA

    ---Purpose: Read & Write tool for FeaSecantCoefficientOfLinearThermalExpansion

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FeaSecantCoefficientOfLinearThermalExpansion from StepFEA

is
    Create returns RWFeaSecantCoefficientOfLinearThermalExpansion from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FeaSecantCoefficientOfLinearThermalExpansion from StepFEA);
	---Purpose: Reads FeaSecantCoefficientOfLinearThermalExpansion

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FeaSecantCoefficientOfLinearThermalExpansion from StepFEA);
	---Purpose: Writes FeaSecantCoefficientOfLinearThermalExpansion

    Share (me; ent : FeaSecantCoefficientOfLinearThermalExpansion from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFeaSecantCoefficientOfLinearThermalExpansion;
