-- File:	MakeParab.cdl
-- Created:	Wed Aug 26 14:31:48 1992
-- Author:	Remi GILET
--		<reg@topsn3>
---Copyright:	 Matra Datavision 1992

class MakeParab from gce inherits Root from gce

    ---Purpose :This class implements the following algorithms used to 
    --          create Parab from gp.
    --  Defines the parabola in the parameterization range  :
    --  ]-infinite, +infinite[
    --  The vertex of the parabola is the "Location" point of the 
    --  local coordinate system (axis placement) of the parabola. 
    --  
    --  The "XDirection" and the "YDirection" of this system define 
    --  the plane of the parabola.
    --  
    --  The "XAxis" of the parabola ("Location", "XDirection") is
    --  the axis of symmetry of the parabola. The Xaxis is oriented 
    --  from the vertex of the parabola to the Focus of the parabola.
    --  
    --  The "YAxis" of the parabola ("Location", "YDirection") is
    --  parallel to the directrix of the parabola.
    --  
    --  The equation of the parabola in the local coordinates system is
    --  Y**2 = (2*P) * X
    --  P is the distance between the focus and the directrix of the 
    --  parabola (called Parameter). 
    --  The focal length F = P/2 is the distance between the vertex 
    --  and the focus of the parabola.
    --          
    --          * Creates a parabola with its local coordinate system "A2"
    --            and it's focal length "Focal".
    --          * Create a parabola with its directrix and its focus point.

uses Pnt   from gp,
     Parab from gp,
     Ax2   from gp,
     Ax1   from gp

raises NotDone from StdFail

is

Create (A2    : Ax2  from gp      ; 
    	Focal : Real from Standard)    returns MakeParab;
    --- Purpose ;
    --  Creates a parabola with its local coordinate system "A2"
    --  and it's focal length "Focal".
    --  The XDirection of A2 defines the axis of symmetry of the 
    --  parabola. The YDirection of A2 is parallel to the directrix
    --  of the parabola. The Location point of A2 is the vertex of
    --  the parabola
    --  The status is "NullFocusLength" if Focal < 0.0


Create (D : Ax1 from gp ; 
    	F : Pnt from gp ) returns MakeParab;
    --- Purpose :
    --  D is the directrix of the parabola and F the focus point.
    --  The symmetry axis (XAxis) of the parabola is normal to the
    --  directrix and pass through the focus point F, but its
    --  location point is the vertex of the parabola.
    --  The YAxis of the parabola is parallel to D and its location
    --  point is the vertex of the parabola. The normal to the plane
    --  of the parabola is the cross product between the XAxis and the
    --  YAxis.

Value(me) returns Parab from gp
    raises NotDone
    is static;
    ---C++: return const&
    ---Purpose: Returns the constructed parabola.
    -- Exceptions StdFail_NotDone if no parabola is constructed.
    
Operator(me) returns Parab from gp
    is static;
    ---C++: return const&
    ---C++: alias "Standard_EXPORT operator gp_Parab() const;"

fields

    TheParab : Parab from gp;
    --The solution from gp.
    
end MakeParab;




