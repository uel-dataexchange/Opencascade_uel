-- File:        SiUnitAndRatioUnit.cdl
-- Created:     Fri Jun 17 11:43:44 1994
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class SiUnitAndRatioUnit from StepBasic inherits SiUnit from StepBasic 

	--- This class is an implementation of EXPRESS
	--  ANDOR Subtype Declaration.
uses

    RatioUnit from StepBasic, 
    DimensionalExponents from StepBasic, 
    SiPrefix from StepBasic, 
    SiUnitName from StepBasic

is

    Create returns mutable SiUnitAndRatioUnit;
	---Purpose: Returns a SiUnitAndRatioUnit

    Init (me: mutable; aDimensions: mutable DimensionalExponents from StepBasic)
    is redefined;

    Init (me: mutable; hasAprefix: Boolean from Standard;
	      	       aPrefix   : SiPrefix from StepBasic;
	      	       aName     : SiUnitName from StepBasic) is redefined;

    -- Specific Methods for Field Data Access --

    SetRatioUnit(me : mutable; aRatioUnit : mutable RatioUnit);
    
    RatioUnit (me) returns mutable RatioUnit;

fields

    ratioUnit: RatioUnit from StepBasic;

end SiUnitAndRatioUnit;
