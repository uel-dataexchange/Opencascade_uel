-- File:	PTopoDS_Shell.cdl
-- Created:	Wed May  5 16:56:49 1993
-- Author:	Remi LEQUETTE
--		<rle@sdsun1>
---Copyright:	 Matra Datavision 1993



class Shell from PTopoDS inherits HShape from PTopoDS

is
    Create returns mutable Shell from PTopoDS;
    ---Level: Internal 

end Shell;
