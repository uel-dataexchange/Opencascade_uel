-- File:        BRepMesh_FastDiscretFace.cdl
-- Created:     Tue Oct 28 14:10:54 2008
-- Author:      
--              <epa@TOSTEX>
---Copyright:    Matra Datavision 2008

private class FastDiscretFace from BRepMesh inherits TShared from MMgt

        ---Purpose: Algorithm  to mesh  a face  with  respect of  the
        --          frontier the deflection  and by option the  shared
        --          components.


uses    Boolean                   from Standard,
        Integer                   from Standard,
        Real                      from Standard,
        Face                      from TopoDS,
        Edge                      from TopoDS,
        Vertex                    from TopoDS,
        Pnt                       from gp,
        Pnt2d                     from gp,
        XY                        from gp,
        HSurface                  from BRepAdaptor,
        Delaun                    from BRepMesh,
        DataStructureOfDelaun     from BRepMesh,
        DataMapOfVertexInteger    from BRepMesh,
        DataMapOfIntegerListOfXY  from BRepMesh,
        DataMapOfShapeReal        from TopTools,
        ListOfVertex              from BRepMesh,
        ClassifierPtr             from BRepMesh,
        Triangle                  from BRepMesh,
        Edge                      from BRepMesh,
        Vertex                    from BRepMesh,
        FaceAttribute             from BRepMesh,
        ListOfInteger             from TColStd,
        BaseAllocator             from BRepMesh,
        DataMapOfIntegerPnt       from BRepMesh,
        IndexedMapOfInteger       from TColStd,
        IndexedMapOfReal          from TColStd,
        DataMapOfShapePairOfPolygon from  BRepMesh,
        Triangulation             from Poly,
        Location                  from TopLoc


is 

        Create (theAngle      : Real    from Standard;
                theWithShare  : Boolean from Standard=Standard_True)
          returns mutable FastDiscretFace from BRepMesh;




        Add  (me       : mutable;
              theFace     : Face from TopoDS;
              theAttrib   : FaceAttribute from BRepMesh;
              theMapDefle : DataMapOfShapeReal from TopTools)
          is static;

      
        Add  (me     : mutable;
              theVert       : Vertex   from TopoDS;
              theFace       : Face     from TopoDS;
              theSFace  : HSurface from BRepAdaptor) is private;
            
        RestoreStructureFromTriangulation
               (me: mutable; 
                theEdge    : Edge          from TopoDS;
                theFace    : Face          from TopoDS;
                theSurf    : HSurface      from BRepAdaptor;
                theTrigu   : Triangulation from Poly;
                theDefEdge : Real          from Standard;
                theLoc     : Location      from TopLoc)
          returns Boolean from Standard is protected;
        
 
        InternalVertices  (me            : mutable;
                           theCaro       : HSurface            from BRepAdaptor;
                           theInternalV  : in out ListOfVertex from BRepMesh;
                           theDefFace    : Real                from Standard;
                           theClassifier : ClassifierPtr       from BRepMesh)
          is static private;


        Control  (me      : mutable;
                  theCaro         : HSurface                from BRepAdaptor;
                  theDefFace      : Real                    from Standard;
                  theInternalV    : in out ListOfVertex     from BRepMesh;
                  theBadTriangles : in out ListOfInteger    from TColStd;
                  theNulTriangles : in out ListOfInteger    from TColStd;
                  theTrigu        : in out Delaun           from BRepMesh;
                  theIsFirst      : Boolean                 from Standard)
          returns Real from Standard is static;

        FindUV (myclass; 
                theV            : Vertex                            from TopoDS; 
                theXY           : Pnt2d                             from gp;
                theIp           : Integer                           from Standard; 
                theSFace        : HSurface                          from BRepAdaptor; 
                theMinDist      : Real                              from  Standard;
                theLocation2dMap: in out DataMapOfIntegerListOfXY   from BRepMesh)
          returns XY from gp;

        AddInShape (me: mutable;
                    theFace   : Face     from TopoDS;
                    theDefFace: Real     from Standard)
          is static private;


-- Output :

        Triangle   (me;
                    theIndex : Integer from Standard)
        ---Purpose: Gives the triangle of <Index>.
        ---C++: return const &
          returns Triangle from BRepMesh
          is static;

        Edge       (me;
                    theIndex : Integer from Standard)
        ---Purpose: Gives the edge of index <Index>.
        ---C++: return const &
          returns Edge from BRepMesh
          is static;


        Vertex     (me;
                    theIndex : Integer from Standard)
          ---Purpose: Gives the vertex of <Index>.
          ---C++: return const &
          returns Vertex from BRepMesh
          is static;

        Pnt        (me;
                    theIndex : Integer from Standard)
          ---Purpose: Gives the location3d of the vertex of <Index>.
          ---C++: return const &
          returns Pnt from gp
          is static;

fields  
        myAngle         : Real                          from Standard;
        myWithShare     : Boolean                       from Standard;
        myVertices      : DataMapOfVertexInteger        from BRepMesh;
        myInternaledges : DataMapOfShapePairOfPolygon   from BRepMesh;
        myNbLocat       : Integer                       from Standard;
        myLocation3d    : DataMapOfIntegerPnt           from BRepMesh;
        myStructure     : DataStructureOfDelaun         from BRepMesh;
        myListver       : ListOfVertex                  from BRepMesh;
        myVemap         : IndexedMapOfInteger           from TColStd;
        myLocation2d    : DataMapOfIntegerListOfXY      from BRepMesh;
        myAttrib        : FaceAttribute                 from BRepMesh;
        myInternalVerticesMode : Boolean                from Standard; --mode to accounting internal vertices 
        myUParam        : IndexedMapOfReal              from TColStd;
        myVParam        : IndexedMapOfReal              from TColStd;
        myAllocator     : BaseAllocator                 from BRepMesh;
 
end FastDiscretFace;
