-- File:	RWStepFEA_RWFeaAxis2Placement3d.cdl
-- Created:	Thu Dec 12 17:51:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFeaAxis2Placement3d from RWStepFEA

    ---Purpose: Read & Write tool for FeaAxis2Placement3d

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FeaAxis2Placement3d from StepFEA

is
    Create returns RWFeaAxis2Placement3d from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FeaAxis2Placement3d from StepFEA);
	---Purpose: Reads FeaAxis2Placement3d

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FeaAxis2Placement3d from StepFEA);
	---Purpose: Writes FeaAxis2Placement3d

    Share (me; ent : FeaAxis2Placement3d from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFeaAxis2Placement3d;
