-- File:        AreaInSet.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWAreaInSet from RWStepVisual

	---Purpose : Read & Write Module for AreaInSet

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     AreaInSet from StepVisual,
     EntityIterator from Interface

is

	Create returns RWAreaInSet;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable AreaInSet from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : AreaInSet from StepVisual);

	Share(me; ent : AreaInSet from StepVisual; iter : in out EntityIterator);

end RWAreaInSet;
