-- File:	IntTools_Compare.cdl
-- Created:	Mon May 22 16:56:20 2000
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2000


class Compare from IntTools 

	---Purpose: Auxiliary class to provide a sorting Roots.     

uses
    Root from IntTools

is
    Create   
    	returns Compare from IntTools;
	---Purpose:
	--- Empty constructor
	---
	 
    Create  (aTol:Real from Standard) 
    	returns Compare from IntTools;
	---Purpose:
	--- Initializes me by tolerance
	---
	 
    IsLower (me; Left, Right: Root from IntTools)
	---Purpose: 
    	--- Returns True if <Left> is lower than <Right>.
	---
    	returns Boolean from Standard;
    
    IsGreater (me; Left, Right: Root from IntTools)
	---Level: Public
	---Purpose: 
    	--- Returns True if <Left> is greater than <Right>.
	---
    	returns Boolean from Standard;

    IsEqual(me; Left, Right: Root from IntTools)
	---Level: Public
	---Purpose: 
    	--- Returns True when <Right> and <Left> are equal.
	---
    	returns Boolean from Standard ;
    	    	

fields
    myTol: Real from Standard; 
     
end Compare;
