-- File:	RWStepAP214_RWAppliedDateAssignment.cdl
-- Created:	Fri Mar 12 11:22:27 1999
-- Author:	data exchange team
--		<det@androx.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999


class RWAppliedDateAssignment from RWStepAP214 

	---Purpose: Read & Write Module for AppliedDateAssignment

uses 
     Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     AppliedDateAssignment from StepAP214,
     EntityIterator from Interface


is
    	Create returns RWAppliedDateAssignment;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable AppliedDateAssignment from StepAP214);

	WriteStep (me; SW : in out StepWriter; ent : AppliedDateAssignment from StepAP214);

	Share(me; ent : AppliedDateAssignment from StepAP214; iter : in out EntityIterator);



end RWAppliedDateAssignment;
