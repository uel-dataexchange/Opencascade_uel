-- File:	StepModel.cdl
-- Created:	Tue Feb 11 16:01:53 1992
-- Author:	Christian CAILLET
--		<cky@phobox>
---Copyright:	 Matra Datavision 1992


class StepModel  from StepData  inherits InterfaceModel

    ---Purpose : Gives access to
    -- - entities in a STEP file,
    -- - the STEP file header.

uses Type, HAsciiString from TCollection,
     Messenger from Message,
     DataMapOfTransientInteger,
     EntityList, EntityIterator, Check

raises NoSuchObject

is

    Create returns mutable StepModel;
    ---Purpose: Creates an empty STEP model with an empty header.
    Reservate (me : mutable; nbent : Integer) is redefined;
    ---Purpose : The standard reservation is completed for the map (id-num)

    Entity (me; num : Integer) returns Transient;
    ---Purpose : returns entity given its rank.
    --           Same as InterfaceEntity, but with a shorter name

    GetFromAnother (me : mutable; other : InterfaceModel);
    ---Purpose : gets header from another Model (uses Header Protocol)

    NewEmptyModel (me) returns mutable InterfaceModel;
    ---Purpose : Returns a New Empty Model, same type as <me>, i.e. StepModel

    	-- --   Header management   -- --

    Header (me) returns EntityIterator;
    ---Purpose : returns Header entities under the form of an iterator

    HasHeaderEntity(me; atype : any Type) returns Boolean;
    ---Purpose : says if a Header entity has a specifed type

    HeaderEntity (me; atype : any Type) returns mutable Transient
    ---Purpose : Returns Header entity with specified type, if there is
    	raises NoSuchObject;
    --           Error if no Header Entity matches <atype>

    ClearHeader (me : mutable);
    ---Purpose : Clears the Header

    AddHeaderEntity (me : mutable; ent : mutable Transient);
    ---Purpose : Adds an Entity to the Header

    VerifyCheck (me; ach : in out Check) is redefined;
    ---Purpose : Specific Check, checks Header Items with HeaderProtocol

    DumpHeader (me; S : Messenger from Message; level : Integer = 0);
    ---Purpose : Dumps the Header, with the Header Protocol of StepData.
    --           If the Header Protocol is not defined, for each Header Entity,
    --           prints its Type. Else sends the Header under the form of
    --           HEADER Section of an Ascii Step File
    --           <level> is not used because Header is not so big


    ClearLabels (me : mutable);
    ---Purpose : erases specific labels, i.e. clears the map (entity-ident)

    SetIdentLabel (me : mutable; ent : Transient; ident : Integer);
    ---Purpose : Attaches an ident to an entity to produce a label
    --           (does nothing if <ent> is not in <me>)

    IdentLabel (me; ent : Transient) returns Integer;
    ---Purpose : returns the label ident attached to an entity, 0 if not in me

    PrintLabel (me; ent : Transient; S : Messenger from Message);
    ---Purpose : Prints label specific to STEP norm for a given entity, i.e.
    --           if a LabelIdent has been recorded, its value with '#', else
    --           the number in the model with '#' and between ()

    StringLabel (me; ent : Transient) returns HAsciiString from TCollection;
    ---Purpose : Returns a string with the label attached to a given entity,
    --           same form as for PrintLabel

fields

    theheader : EntityList;
    theidnums : DataMapOfTransientInteger;

end StepModel;
