
-- File:	Graphic2d_Buffer.cdl
-- Created:	Mercredi 15 fevrier 1995
-- Authors:	CAL, GG
--
---Copyright:	Matra Datavision 1995

class Buffer from Graphic2d inherits TShared from MMgt

    	---Purpose: This class constructs a 2D graphic buffer in a view.   It
    	-- manages a set of graphic objects and/or primitives.
    	-- To draw the buffer, the following elements are required:
    	-- -   the override color
    	-- -   the font
    	-- -   a solid line type
    	-- -   thickness of 1 pixel.
    	-- With this category , the user can drag the geometry
    	-- stored in the buffer without changing the fixed
    	-- background.   This mechanism is reserved for the
    	-- special driver Aspect_WindowDriver:   if no other
    	-- driver has been defined, nothing will be drawn.   Both
    	-- this driver and view mapping are used to draw the buffer.
    	-- Warning
    	-- -   This class manages dragging only.   It does not
    	--   manage "sketching" or "rubberbanding".   For example:
    	--   -   There is no empty constructor for this
    	--    primitive.   Therefore we must create a primitive
    	--    in a dummy object simply to add this primitive to the buffer.
    	--   -   There is no Buffer->Add (anArrayOfPoints)
    	--    method.   Therefor it is not possible to add
    	--    shapes to the buffer.
    	--   -   There are no Polyline->ChangeApoint () nor
    	--    Circle->ChangeRadius () methods.   Therefore
    	--    we must call the primitive's destructor to modify
    	--    the definition of one primitive in a buffer.
    	-- -   The Graphic2d_Image class is a primitive.   For
    	--   this class, we replace the definition of the image
    	--   with a rectangle with the same size and the same position.
    	-- -   You can add or remove primitives to the buffer
    	--   after creating and displaying it again.
        
        
        
uses
	PlaneAngle		from Quantity,
	Factor			from Quantity,
	Length			from Quantity,

	View			from Graphic2d,
	Drawer			from Graphic2d,
	ViewPtr			from Graphic2d,
	Primitive		from Graphic2d,
	SequenceOfPrimitives	from Graphic2d,
	GraphicObject		from Graphic2d,
	SequenceOfGraphicObject from Graphic2d,
	ViewMapping 		from Graphic2d,
	WindowDriver		from Aspect,
	TypeOfDrawMode		from Aspect

is
	-------------------------
	-- Category: Constructors
	-------------------------

	Create (aView: View from Graphic2d;
		aPivotX, aPivotY: Length from Quantity;
		aWidthIndex: Integer from Standard = 0;
		aColorIndex: Integer from Standard = 0;
		aFontIndex: Integer from Standard = 0;
		aDrawMode: TypeOfDrawMode from Aspect = Aspect_TODM_REPLACE)
	returns mutable Buffer from Graphic2d;
	---Purpose:	Creates an empty graphic buffer in the view <aView>.
	--		A graphic buffer manages a set of graphic objects
	--		and/or primitives.
	--		A buffer color and font index can be defined,
	--		in place of the default overrideColor or systemFont.
	--		When the drawmode is REPLACE the buffer is drawn with
	--		the right color and background drawing is used for 
	--		restoring it at Erase() time.
	--		When the drawmode is XOR the buffer is drawn or erase
	--		with an optimal color depending of the background color
	--		but some side effects can appears depending of
	--		background drawing pixels values.
	---Category:	Constructors

	------------------------
	-- Category: Destructors
	------------------------

	Destroy (me: mutable)
	is static;
	---Level:	Public
	---Purpose:	Deletes the graphic buffer <me>.
	---C++:		alias ~
	---Category:	Destructors

	---------------------------------------------------------
	-- Category: Methods to manage the contents of the buffer
	---------------------------------------------------------

	Add (me: mutable; anObject: GraphicObject from Graphic2d)
	is static;
	---Level:	Public
	---Purpose:	Adds the graphic object <anObject> in the graphic
	--		buffer <me>.
	---Category:	Methods to manage the contents of the buffer

	Add (me: mutable; aPrimitive: Primitive from Graphic2d)
	is static;
	---Level:	Public
	---Purpose:	Adds the primitive <aPrimitive> in the graphic
	--		buffer <me>.
	---Category:	Methods to manage the contents of the buffer

	Remove (me: mutable; anObject: GraphicObject from Graphic2d)
	is static;
	---Level:       Public
        ---Purpose:     Removes the object <anObject> from the graphic
        --              buffer <me>.
        ---Category:    Methods to manage the contents of the buffer

        Remove (me: mutable; aPrimitive: Primitive from Graphic2d)
        is static;
        ---Level:       Public
        ---Purpose:     Removes the primitive <aPrimitive> from the graphic
        --              buffer <me>.
        ---Category:    Methods to manage the contents of the buffer

	Clear (me: mutable)
	is static;
	---Level:	Public
	---Purpose:	Clears the graphic buffer <me>.
	--		Removes all the primitives from the graphic buffer <me>.
	---Category:	Methods to manage the contents of the buffer
--
	---------------------------------------------------------
	-- Category: Methods to manage the attributes of the buffer
	---------------------------------------------------------

	SetAttrib(me : mutable;
		aWidthIndex: Integer from Standard;
		aColorIndex: Integer from Standard;
		aFontIndex: Integer from Standard;
		aDrawMode: TypeOfDrawMode from Aspect) is static;
	---Level:	Public
	---Purpose:	Updates the default buffer color with a new
	--		color index defines in the user ColorMap.
	--         	Update the default buffer font with a new
	--		font index defines in the user FontMap.
	--		Update the default buffer drawmode with
	--		REPLACE or XOR .
	--		You can specify the width index
	--		- -1 draw all lines with the largest width
	--		  defined in the buffer <me>
	--		- 0 draw all lines with the default width
	--		  defined in the driver (1 pixel)
	--		- draw all lines with the specified width
	--		  <aWidthIndex>
	--		You can specify the color index
	--		- -1 draw all primitives with the color of
	--		  the first primitive color defined in the buffer.
	--		- 0 draw all primitives with the default color.
	--		You can specify the font index
	--		- -1 draw all text primitives with the font of
	--		  the first primitive text defined in the buffer.
	--		- 0 draw all text primitives with the default font.
	--  Warning:	The buffer is redisplayed again if it was posted.
	---Category:	Methods to manage the attributes of the buffer

	SetPivot(me : mutable;
		aPivotX, aPivotY: Length from Quantity)
	is static;
	---Level:	Public
	---Purpose:	Updates the buffer pivot position.
	--  Warning:	The buffer is redisplayed again if it was posted.
	---Category:	Methods to manage the position of the buffer

	SetPivot(me : mutable)
	is static;
	---Level:	Public
	---Purpose:	Updates the buffer pivot position with the actual position.
	---Category:	Methods to manage the position of the buffer

--
	---------------------------------------------------------
	-- Category: Methods to manage the position of the buffer
	---------------------------------------------------------

	Move (me: mutable;
		aDeltaX,aDeltaY: Length from Quantity)
	is static;
	---Level:	Public
	---Purpose:	Moves the graphic buffer <me> at the specified
	--		position. The new position of the buffer is :
	--		(<aPivotX> + <aDeltaX>, <aPivotY> + <aDeltaY>)
	---Category:	Methods to manage the position of the buffer

	Rotate (me: mutable;
		anAngle: PlaneAngle from Quantity)
	is static;
	---Level:	Public
	---Purpose:	Rotates the graphic buffer <me> with the specified
	--		absolute counter clockwise angle from the pivot X axis.
	---Category:	Methods to manage the position of the buffer

	Scale (me: mutable;
		aFactor: Factor from Quantity)
	is static;
	---Level:	Public
	---Purpose:	Scales the graphic buffer <me> with the specified
	--		absolute scale factor from the pivot point.
	---Category:	Methods to manage the position of the buffer

	----------------------------
	-- Category: Inquire methods
	----------------------------

	View (me)
	returns mutable View from Graphic2d is static;
	---Level:	Public
	---Purpose:	Returns the view which manages the graphic buffer <me>.
	---Category:	Inquire methods

	IsEmpty (me)
	returns Boolean from Standard
	is static;
	---Level:	Public
	---Purpose:	Returns Standard_True if the graphic buffer <me>
	--		is empty, Standard_False if not.
	---Category:	Inquire methods

	IsIn (me; aPrimitive: Primitive from Graphic2d)
	returns Boolean from Standard
	is static;
	---Level:	Public
	---Purpose:	Returns Standard_True if the primitive <aPrimitive>
	--		is in the graphic buffer <me>, Standard_False if not.
	---Category:	Inquire methods

	IsIn (me; anObject: GraphicObject from Graphic2d)
	returns Boolean from Standard
	is static;
	---Level:	Public
	---Purpose:	Returns Standard_True if the graphic object <anObject>
	--		is in the graphic buffer <me>, Standard_False if not.
	---Category:	Inquire methods

	---------------------------------------------
	-- Category: Methods to manage the visibility
	---------------------------------------------

	Post (me: mutable)
	is static;
	---Level:	Public
	---Purpose:	Post the graphic buffer in the current View driver
	-- and display it.
	--  Warning: The view driver must be defined and of type WindowDriver
	-- or nothing is drawn .
	---Category:	Methods to manage the visibility

	Post (me: mutable;
                aDriver: WindowDriver from Aspect;
                aViewMapping: ViewMapping from Graphic2d;
                aXPosition, aYPosition: Real from Standard;
                aScale: Real from Standard)
	is static;
	---Level:	Public
	---Purpose:	Post the graphic buffer in a View driver and display it.
	---Category:	Methods to manage the visibility

	UnPost (me: mutable)
	is static;
	---Level:	Public
	---Purpose:	Unpost the graphic buffer from the view and erase it.
	---Category:	Methods to manage the visibility

	IsPosted (me)
	returns Boolean from Standard
	is static;
	---Level:	Public
	---Purpose:	Returns Standard_True if the graphic buffer <me>
	--		is posted in the view, Standard_False if not.
	---Category:	Methods to manage the visibility

	IsPosted (me;
                aDriver: WindowDriver from Aspect)
	returns Boolean from Standard
	is static private;
	---Level:	Public
	---Purpose:	Returns Standard_True if the graphic buffer <me>
	--		is posted in the view with the driver <aDriver>, 
	--		Standard_False if not.
	---Category:	Private methods

	-------------------------------------------------------------
	-- Category: Inquiries to retrieve the position of the buffer
	-------------------------------------------------------------

	Angle (me)
	returns PlaneAngle from Quantity is static;
	---Level:	Public
	---Purpose:	Returns the value of the rotation angle of the
	--		graphic buffer <me>.
	---Category:	Inquire methods

	Scale (me)
	returns Factor from Quantity is static;
	---Level:	Public
	---Purpose:	Returns the value of the scale factor of the
	--		graphic buffer <me>.
	---Category:	Inquire methods

	Xpivot (me)
	returns Length from Quantity is static;
	---Level:	Public
	---Purpose:	Returns the actual value of the X pivot point.
	--		of the graphic buffer <me>.
	---Category:	Inquire methods

	Ypivot (me)
	returns  Length from Quantity is static;
	---Level:	Public
	---Purpose:	Returns the actual value of the Y pivot point.
	--		of the graphic buffer <me>.
	---Category:	Inquire methods

	----------------------------
	-- Category: Private methods
	----------------------------

	Draw (me : mutable) is static private;
	---Level:	Internal
	---Purpose:	Update the internal buffer with new primitives
	--		if any and draw it at screen.
	---Category:	Private methods

	Erase (me : mutable) is static private;
	---Level:	Internal
	---Purpose:	Erase the internal buffer from the screen.
	---Category:	Private methods

	ReLoad (me : mutable; 
		ResetPosition: Boolean from Standard = Standard_True) 
		is static private;
	---Level:	Internal
	---Purpose:	Erase and Reload the internal graphic buffer before
	--		drawing to the current drawer.
	--		Keep the actual position if <ResetPosition> is FALSE.
	---Category:	Private methods

	MaxWidth (me; theWidth: out Length from Quantity;
		      theIndex: out Integer from Standard)
	returns Boolean from Standard is static private;
	---Level:	Internal
	---Purpose:	Returns Standard_True if the buffer contains
	--		lines and the maximum width of the lines in the
	--		buffer <me>
	---Category:	Private methods

fields
	myBufferId:		Integer from Standard;
	myBufferIsPosted:	Boolean from Standard;
	myDriver:		WindowDriver from Aspect;
	myPivotX:		ShortReal from Standard;
	myPivotY:		ShortReal from Standard;
	myWidthIndex:		Integer from Standard;
	myColorIndex:		Integer from Standard;
	myFontIndex:		Integer from Standard;
	myDrawMode:		TypeOfDrawMode from Aspect;
	myPView:		ViewPtr from Graphic2d;
	myPrimitives:		SequenceOfPrimitives from Graphic2d;
	myObjects:		SequenceOfGraphicObject from Graphic2d;

friends

	class View from Graphic2d

end Buffer from Graphic2d;
