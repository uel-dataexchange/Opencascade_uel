-- File:	BinTools_SurfaceSet.cdl
-- Created:	Thu May 20 14:33:11 2004
-- Author:	Sergey ZARITCHNY <szy@opencascade.com>
-- Copyright:	Open CasCade S.A. 2004 


class SurfaceSet from BinTools  

	---Purpose: Stores a set of Surfaces from Geom in binary format.

uses
    Surface from Geom,
    IndexedMapOfTransient from TColStd
    
raises
    OutOfRange from Standard

is

    Create returns SurfaceSet from BinTools;
	---Purpose: Returns an empty set of Surfaces.
	
    Clear(me : in out)
	---Purpose: Clears the content of the set.
    is static;
	
    Add(me : in out; S : Surface from Geom) returns Integer
	---Purpose: Incorporate a new Surface in the  set and returns
	--          its index.
    is static;
    
    Surface(me; I : Integer) returns Surface from Geom
	---Purpose: Returns the Surface of index <I>.
    raises
    	OutOfRange from Standard
    is static;

    Index(me; S : Surface from Geom) returns Integer
	---Purpose: Returns the index of <L>.
    is static;
    	
    Write(me; OS : in out OStream)
	---Purpose: Writes the content of  me  on the stream <OS> in 
	--          binary format that can be read back by Read.
    is static;
	
    Read(me : in out; IS : in out IStream)
	---Purpose: Reads the content of me from the  stream  <IS>. me
	--          is first cleared.
	--          
    is static;
	
    --
    -- 	class methods to write an read surfaces
    -- 	
    
    WriteSurface(myclass; S  : Surface from Geom;
    	    	    	  OS : in out OStream);
	---Purpose: Dumps the surface on the stream in binary
	--          format that can be read back.
	
    ReadSurface(myclass; IS : in out IStream;
    	    	         S  : in out Surface from Geom)
    returns IStream;
	---Purpose: Reads the surface  from  the stream.  The  surface  is
	--          assumed   to have  been  written  with  the Write
	--          method.
	--          
	---C++: return &
	
fields

    myMap : IndexedMapOfTransient from TColStd;

end SurfaceSet;
