-- File:	RWStepElement_RWVolume3dElementDescriptor.cdl
-- Created:	Thu Dec 12 17:29:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWVolume3dElementDescriptor from RWStepElement

    ---Purpose: Read & Write tool for Volume3dElementDescriptor

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    Volume3dElementDescriptor from StepElement

is
    Create returns RWVolume3dElementDescriptor from RWStepElement;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : Volume3dElementDescriptor from StepElement);
	---Purpose: Reads Volume3dElementDescriptor

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: Volume3dElementDescriptor from StepElement);
	---Purpose: Writes Volume3dElementDescriptor

    Share (me; ent : Volume3dElementDescriptor from StepElement;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWVolume3dElementDescriptor;
