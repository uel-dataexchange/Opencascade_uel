-- File:	IGESAppli_ToolNodalResults.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolNodalResults  from IGESAppli

    ---Purpose : Tool to work on a NodalResults. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses NodalResults from IGESAppli,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolNodalResults;
    ---Purpose : Returns a ToolNodalResults, ready to work


    ReadOwnParams (me; ent : mutable NodalResults;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : NodalResults;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : NodalResults;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a NodalResults <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : NodalResults) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : NodalResults;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : NodalResults; entto : mutable NodalResults;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : NodalResults;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolNodalResults;
