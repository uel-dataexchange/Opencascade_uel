-- File:        BoundedCurve.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWBoundedCurve from RWStepGeom

	---Purpose : Read & Write Module for BoundedCurve

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     BoundedCurve from StepGeom

is

	Create returns RWBoundedCurve;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable BoundedCurve from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : BoundedCurve from StepGeom);

end RWBoundedCurve;
