-- File:        AutoDesignActualDateAndTimeAssignment.cdl
-- Created:     Fri Dec  1 11:11:13 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class AutoDesignActualDateAndTimeAssignment from StepAP214 

inherits DateAndTimeAssignment from StepBasic 

uses

	HArray1OfAutoDesignDateAndTimeItem from StepAP214, 
	AutoDesignDateAndTimeItem from StepAP214, 
	DateAndTime from StepBasic, 
	DateTimeRole from StepBasic
is

	Create returns mutable AutoDesignActualDateAndTimeAssignment;
	---Purpose: Returns a AutoDesignActualDateAndTimeAssignment


	Init (me : mutable;
	      aAssignedDateAndTime : mutable DateAndTime from StepBasic;
	      aRole : mutable DateTimeRole from StepBasic) is redefined;

	Init (me : mutable;
	      aAssignedDateAndTime : mutable DateAndTime from StepBasic;
	      aRole : mutable DateTimeRole from StepBasic;
	      aItems : mutable HArray1OfAutoDesignDateAndTimeItem from StepAP214) is virtual;

	-- Specific Methods for Field Data Access --

	SetItems(me : mutable; aItems : mutable HArray1OfAutoDesignDateAndTimeItem);
	Items (me) returns mutable HArray1OfAutoDesignDateAndTimeItem;
	ItemsValue (me; num : Integer) returns AutoDesignDateAndTimeItem;
	NbItems (me) returns Integer;

fields

	items : HArray1OfAutoDesignDateAndTimeItem from StepAP214; -- a SelectType

end AutoDesignActualDateAndTimeAssignment;
