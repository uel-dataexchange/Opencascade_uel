-- File:	RWStepFEA_RWFeaParametricPoint.cdl
-- Created:	Thu Dec 12 17:51:06 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFeaParametricPoint from RWStepFEA

    ---Purpose: Read & Write tool for FeaParametricPoint

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FeaParametricPoint from StepFEA

is
    Create returns RWFeaParametricPoint from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FeaParametricPoint from StepFEA);
	---Purpose: Reads FeaParametricPoint

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FeaParametricPoint from StepFEA);
	---Purpose: Writes FeaParametricPoint

    Share (me; ent : FeaParametricPoint from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFeaParametricPoint;
