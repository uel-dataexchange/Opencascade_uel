-- File:	IGESDimen_ToolBasicDimension.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolBasicDimension  from IGESDimen

    ---Purpose : Tool to work on a BasicDimension. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses BasicDimension from IGESDimen,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolBasicDimension;
    ---Purpose : Returns a ToolBasicDimension, ready to work


    ReadOwnParams (me; ent : mutable BasicDimension;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : BasicDimension;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : BasicDimension;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a BasicDimension <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable BasicDimension) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a BasicDimension
    --           (NbPropertyValues forced to 8)

    DirChecker (me; ent : BasicDimension) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : BasicDimension;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : BasicDimension; entto : mutable BasicDimension;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : BasicDimension;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolBasicDimension;
