-- File:	RWStepRepr_RWShapeAspectTransition.cdl
-- Created:	Tue Apr 18 16:42:58 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWShapeAspectTransition from RWStepRepr

    ---Purpose: Read & Write tool for ShapeAspectTransition

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ShapeAspectTransition from StepRepr

is
    Create returns RWShapeAspectTransition from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ShapeAspectTransition from StepRepr);
	---Purpose: Reads ShapeAspectTransition

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ShapeAspectTransition from StepRepr);
	---Purpose: Writes ShapeAspectTransition

    Share (me; ent : ShapeAspectTransition from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWShapeAspectTransition;
