-- File:	StepToGeom_MakeSurfaceOfLinearExtrusion.cdl
-- Created:	Mon Jun 14 16:16:49 1993
-- Author:	Martine LANGLOIS
---Copyright:	 Matra Datavision 1993

class MakeSurfaceOfLinearExtrusion from StepToGeom

    ---Purpose: This class implements the mapping between class
    --          SurfaceOfLinearExtrusion from StepGeom which describes a
    --          surface_of_linear_extrusion from Prostep and 
    --          SurfaceOfLinearExtrusion from Geom.

uses SurfaceOfLinearExtrusion from Geom,
     SurfaceOfLinearExtrusion from StepGeom

is 

    Convert ( myclass; SS : SurfaceOfLinearExtrusion from StepGeom;
                       CS : out SurfaceOfLinearExtrusion from Geom )
    returns Boolean from Standard;

end MakeSurfaceOfLinearExtrusion;
