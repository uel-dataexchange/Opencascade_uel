-- File:        GeometricallyBoundedWireframeShapeRepresentation.cdl
-- Created:     Fri Dec  1 11:11:21 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class GeometricallyBoundedWireframeShapeRepresentation from StepShape 

inherits ShapeRepresentation from StepShape 

uses

	HAsciiString from TCollection, 
	HArray1OfRepresentationItem from StepRepr,
	RepresentationContext from StepRepr
is

	Create returns mutable GeometricallyBoundedWireframeShapeRepresentation;
	---Purpose: Returns a GeometricallyBoundedWireframeShapeRepresentation


end GeometricallyBoundedWireframeShapeRepresentation;
