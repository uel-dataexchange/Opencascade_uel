-- File:	STEPEdit.cdl
-- Created:	Wed Jul 29 11:56:51 1998
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1998


package STEPEdit

    ---Purpose : Provides tools to exploit and edit a set of STEP data :
    --           editors, selections ..

uses Standard, TCollection,
     Interface, IFSelect, StepData

is

    class EditContext;
    -- This class is for global context : ApplicationContext,
    --   ProductRelatedProductCategory

    class EditSDR;
    -- This class allows to edit product data for a SDR


    	--  Some useful operators
    	--  They are not classes, they are just based on general tools

    Protocol returns Protocol from Interface;
    ---Purpose : Returns a Protocol fit for STEP (creates the first time)

    NewModel returns StepModel from StepData;
    ---Purpose : Returns a new empty StepModel fit for STEP
    --           i.e. with its header determined from Protocol

    SignType returns Signature from IFSelect;
    ---Purpose : Returns a SignType fit for STEP (creates the first time)

    NewSelectSDR returns SelectSignature from IFSelect;
    ---Purpose : Creates a Selection for ShapeDefinitionRepresentation
    --           By default searches among root entities

    NewSelectPlacedItem returns SelectSignature from IFSelect;
    ---Purpose : Creates a Selection for Placed Items, i.e. MappedItem or
    --           ContextDependentShapeRepresentation, which itself refers to a
    --           RepresentationRelationship with possible subtypes (Shape...
    --           and/or ...WithTransformation)
    --           By default in the whole StepModel

    NewSelectShapeRepr returns SelectSignature from IFSelect;
    ---Purpose : Creates a Selection for ShapeRepresentation and its sub-types,
    --           plus ContextDependentShapeRepresentation (which is not a
    --           sub-type of ShapeRepresentation)
    --           By default in the whole StepModel

end STEPEdit;
