-- File:	RWStepRepr_RWConfigurationItem.cdl
-- Created:	Fri Nov 26 16:26:37 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWConfigurationItem from RWStepRepr

    ---Purpose: Read & Write tool for ConfigurationItem

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ConfigurationItem from StepRepr

is
    Create returns RWConfigurationItem from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ConfigurationItem from StepRepr);
	---Purpose: Reads ConfigurationItem

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ConfigurationItem from StepRepr);
	---Purpose: Writes ConfigurationItem

    Share (me; ent : ConfigurationItem from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWConfigurationItem;
