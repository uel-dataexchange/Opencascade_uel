-- File:	TDocStd_Owner.cdl
-- Created:	Mon Jul 12 08:39:13 1999
-- Author:	Denis PASCAL
--		<dp@dingox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1999



private class Owner from TDocStd inherits Attribute from TDF

	---Purpose: 

uses Attribute from TDF,
     GUID      from Standard, 
     RelocationTable from TDF, 
     Data      from TDF,
     Label     from TDF,
     Document  from TDocStd

is 

    ---Purpose: class methods
    --          =============

    GetID (myclass)   
    	---C++: return const &  
    returns GUID from Standard;

    SetDocument (myclass; indata : Data from TDF; doc : Document from TDocStd);
    
    GetDocument (myclass; ofdata : Data from TDF)
    returns Document from TDocStd;

    ---Purpose: Owner methods
    --          ===============
    
    Create
    returns mutable Owner from TDocStd;  
    
    SetDocument (me : mutable; document : Document from TDocStd);    

    GetDocument (me)
    returns Document from TDocStd;
    
    ---Category: methodes de TDF_Attribute
    --           =========================
    
    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; Into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

    Dump(me; anOS : in out OStream from Standard)
    	returns OStream from Standard
    	is redefined;
	---C++: return &

fields

    myDocument : Document from TDocStd;

end Owner;
