-- File:	RWStepFEA_RWCurveElementEndOffset.cdl
-- Created:	Thu Dec 12 17:51:03 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWCurveElementEndOffset from RWStepFEA

    ---Purpose: Read & Write tool for CurveElementEndOffset

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    CurveElementEndOffset from StepFEA

is
    Create returns RWCurveElementEndOffset from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : CurveElementEndOffset from StepFEA);
	---Purpose: Reads CurveElementEndOffset

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: CurveElementEndOffset from StepFEA);
	---Purpose: Writes CurveElementEndOffset

    Share (me; ent : CurveElementEndOffset from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWCurveElementEndOffset;
