-- File:	IGESDimen_ToolNewDimensionedGeometry.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolNewDimensionedGeometry  from IGESDimen

    ---Purpose : Tool to work on a NewDimensionedGeometry. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses NewDimensionedGeometry from IGESDimen,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolNewDimensionedGeometry;
    ---Purpose : Returns a ToolNewDimensionedGeometry, ready to work


    ReadOwnParams (me; ent : mutable NewDimensionedGeometry;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : NewDimensionedGeometry;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : NewDimensionedGeometry;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a NewDimensionedGeometry <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable NewDimensionedGeometry) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a NewDimensionedGeometry
    --           (NbDimensions forced to 1, Transf Nullified in D.E.)

    DirChecker (me; ent : NewDimensionedGeometry) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : NewDimensionedGeometry;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : NewDimensionedGeometry; entto : mutable NewDimensionedGeometry;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : NewDimensionedGeometry;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolNewDimensionedGeometry;
