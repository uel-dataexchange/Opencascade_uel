-- File:	StepShape_ConnectedFaceSubSet.cdl
-- Created:	Fri Jan  4 17:42:43 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class ConnectedFaceSubSet from StepShape
inherits ConnectedFaceSet from StepShape

    ---Purpose: Representation of STEP entity ConnectedFaceSubSet

uses
    HAsciiString from TCollection,
    HArray1OfFace from StepShape,
    ConnectedFaceSet from StepShape

is
    Create returns ConnectedFaceSubSet from StepShape;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aConnectedFaceSet_CfsFaces: HArray1OfFace from StepShape;
                       aParentFaceSet: ConnectedFaceSet from StepShape);
	---Purpose: Initialize all fields (own and inherited)

    ParentFaceSet (me) returns ConnectedFaceSet from StepShape;
	---Purpose: Returns field ParentFaceSet
    SetParentFaceSet (me: mutable; ParentFaceSet: ConnectedFaceSet from StepShape);
	---Purpose: Set field ParentFaceSet

fields
    theParentFaceSet: ConnectedFaceSet from StepShape;

end ConnectedFaceSubSet;
