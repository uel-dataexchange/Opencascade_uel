-- File:	RWStepFEA_RWSurface3dElementRepresentation.cdl
-- Created:	Thu Dec 12 17:51:07 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWSurface3dElementRepresentation from RWStepFEA

    ---Purpose: Read & Write tool for Surface3dElementRepresentation

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    Surface3dElementRepresentation from StepFEA

is
    Create returns RWSurface3dElementRepresentation from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : Surface3dElementRepresentation from StepFEA);
	---Purpose: Reads Surface3dElementRepresentation

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: Surface3dElementRepresentation from StepFEA);
	---Purpose: Writes Surface3dElementRepresentation

    Share (me; ent : Surface3dElementRepresentation from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWSurface3dElementRepresentation;
