-- File:	STEPControl_Writer.cdl
-- Created:	Mon Jul  8 16:13:44 1996
-- Author:	Christian CAILLET
--		<cky@anion.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996


class Writer from STEPControl

    	---Purpose : This class creates and writes
    	-- STEP files from Open CASCADE models. A STEP file can be
    	-- written to an existing STEP file or to a new one.
    	-- Translation can be performed in one or several operations. Each
    	-- translation operation outputs a distinct root entity in the STEP file.

uses

    CString,
    StepModel from StepData, WorkSession from XSControl,
    ReturnStatus from IFSelect,
    Shape from TopoDS,
    StepModelType from STEPControl

is

    Create returns Writer;
    ---Purpose : Creates a Writer from scratch

    Create (WS : mutable WorkSession from XSControl;
    	    	 scratch : Boolean = Standard_True) returns Writer;
    ---Purpose : Creates a Writer from an already existing Session
    --           If <scratch> is True (D), clears already recorded data

    SetTolerance (me : in out; Tol : Real);
    ---Purpose : Sets a length-measure value that
    --           will be written to uncertainty-measure-with-unit
    --           when the next shape is translated.

    UnsetTolerance (me : in out);
    ---Purpose : Unsets the tolerance formerly forced by SetTolerance

    SetWS (me : in out; WS : mutable WorkSession from XSControl;
    	    	 scratch : Boolean = Standard_True);
    ---Purpose : Sets a specific session to <me>

    WS (me) returns WorkSession from XSControl;
    ---Purpose : Returns the session used in <me>

    Model (me : in out; newone : Boolean = Standard_False) returns StepModel;
    ---Purpose : Returns the produced model. Produces a new one if not yet done
    --           or if <newone> is True
    --           This method allows for instance to edit product or header
    --           data before writing.

    Transfer (me : in out; sh : Shape from TopoDS;
    	    	    	   mode : StepModelType from STEPControl;
    	    	    	   compgraph : Boolean = Standard_True)
    	returns ReturnStatus;
    	---Purpose : Translates shape sh to a STEP
    	-- entity. mode defines the STEP entity type to be output:
    	-- - STEPControlStd_AsIs translates a shape to its highest possible
    	--   STEP representation.
    	-- - STEPControlStd_ManifoldSolidBrep translates a shape to a STEP
    	--   manifold_solid_brep or brep_with_voids entity.
    	-- - STEPControlStd_FacetedBrep translates a shape into a STEP
    	--   faceted_brep entity.
    	-- - STEPControlStd_ShellBasedSurfaceModel translates a shape into a STEP
    	--   shell_based_surface_model entity.
    	-- - STEPControlStd_GeometricCurveSet translates a shape into a STEP
    	--   geometric_curve_set entity.
  

    Write (me : in out; filename : CString) returns ReturnStatus;
    	---Purpose : Writes a STEP model in the file identified by filename.

    PrintStatsTransfer (me; what : Integer; mode : Integer = 0);
    	---Purpose :  Displays the statistics for the
    	-- last translation. what defines the kind of statistics that are displayed:
    	-- - 0 gives general statistics   (number of translated roots,
    	--   number of warnings, number of   fail messages),
    	-- - 1 gives root results,
    	-- - 2 gives statistics for all checked entities,
    	-- - 3 gives the list of translated entities,
    	-- - 4 gives warning and fail messages,
    	-- - 5 gives fail messages only.
    	--   mode is used according to the use of what. If what is 0, mode is
    	-- ignored. If what is 1, 2 or 3, mode defines the following:
    	-- - 0 lists the numbers of STEP entities in a STEP model,
    	-- - 1 gives the number, identifier, type and result type for each
    	--   STEP entity and/or its status (fail, warning, etc.),
    	-- - 2 gives maximum information for each STEP entity (i.e. checks),
    	-- - 3 gives the number of entities by the type of a STEP entity,
    	-- - 4 gives the number of of STEP entities per result type and/or status,
    	-- - 5 gives the number of pairs (STEP or result type and status),
    	-- - 6 gives the number of pairs (STEP or result type and status)
    	--   AND the list of entity numbers in the STEP model.

fields

    thesession : WorkSession from XSControl;

end Writer;
