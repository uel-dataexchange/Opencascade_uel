-- File:	BinXCAFDrivers_DocumentStorageDriver.cdl
-- Created:	Mon Apr 18 17:07:18 2005
-- Author:	Eugeny NAPALKOV <eugeny.napalkov@opencascade.com>
-- Copyright:	Open CasCade S.A. 2005

class DocumentStorageDriver from BinXCAFDrivers inherits DocumentStorageDriver from BinDrivers

uses
    MessageDriver    from CDM,
    ADriverTable     from BinMDF
is

    Create returns mutable DocumentStorageDriver from BinXCAFDrivers;
	---Purpose: Constructor


    AttributeDrivers  (me : mutable; theMsgDriver: MessageDriver from CDM)
	returns ADriverTable from BinMDF
	is redefined virtual;

end DocumentStorageDriver;

