-- File:	StepBasic_MeasureValueMember.cdl
-- Created:	Fri Mar 28 10:57:37 1997
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


class MeasureValueMember  from StepBasic    inherits  SelectReal  from StepData

    ---Purpose : for Select MeasureValue, i.e. :
    --         length_measure,time_measure,plane_angle_measure,
    --         solid_angle_measure,ratio_measure,parameter_value,
    --         context_dependent_measure,positive_length_measure,
    --         positive_plane_angle_measure,positive_ratio_measure,
    --	       area_measure,volume_measure

uses CString

is

    Create returns mutable MeasureValueMember;
    -- starts as case null (no name)

    HasName (me) returns Boolean  is redefined;
    -- returns True is case not null

    Name    (me) returns CString  is redefined;
    --  returns a name according to the case
    --  0 -> void
    --  1 -> LENGTH_MEASURE
    --  2 -> TIME_MEASURE
    --  3 -> PLANE_ANGLE_MEASURE
    --  4 -> SOLID_ANGLE_MEASURE
    --  5 -> RATIO_MEASURE
    --  6 -> PARAMETER_VALUE
    --  7 -> CONTEXT_DEPENDANT_MEASURE
    --  8 -> POSITIVE_LENGTH_MEASURE
    --  9 -> POSITIVE_PLANE_ANGLE_MEASURE
    --  10 -> POSITIVE_RATIO_MEASURE
    --  11 -> AREA_MEASURE
    --  12 ->VOLUME_MEASURE
    --  13 ->MASS_MEASURE
    --  14 ->THERMODYNAMIC_TEMPERATURE_MEASURE
    
    SetName (me : mutable; name : CString)  returns Boolean  is redefined;
    -- checks for one of the names above, and sets the case number
    -- accepts a void name (case 0)

fields

    thecase : Integer;

end MeasureValueMember;
