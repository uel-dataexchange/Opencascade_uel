-- File:	BinMXCAFDoc_DocumentToolDriver.cdl
-- Created:	Tue May 17 12:26:47 2005
-- Author:	Eugeny NAPALKOV <eugeny.napalkov@opencascade.com>
-- Copyright:	Open CasCade S.A. 2005

class DocumentToolDriver from BinMXCAFDoc inherits ADriver from BinMDF

uses
    MessageDriver    from CDM,
    SRelocationTable from BinObjMgt,
    RRelocationTable from BinObjMgt,
    Persistent       from BinObjMgt,
    Attribute        from TDF

is
    Create (theMsgDriver:MessageDriver from CDM)
    returns mutable DocumentToolDriver from BinMXCAFDoc;

    NewEmpty (me)  returns mutable Attribute from TDF
    is redefined;

    Paste(me; theSource     : Persistent from BinObjMgt;
              theTarget     : mutable Attribute from TDF;
              theRelocTable : out RRelocationTable from BinObjMgt)
    returns Boolean from Standard is redefined;

    Paste(me; theSource     : Attribute from TDF;
              theTarget     : in out Persistent from BinObjMgt;
              theRelocTable : out SRelocationTable from BinObjMgt)
    is redefined;

end;

