-- File:        ProductDefinitionFormationWithSpecifiedSource.cdl
-- Created:     Fri Dec  1 11:11:26 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class ProductDefinitionFormationWithSpecifiedSource from StepBasic 

inherits ProductDefinitionFormation from StepBasic 

uses

	Source from StepBasic, 
	HAsciiString from TCollection, 
	Product from StepBasic
is

	Create returns mutable ProductDefinitionFormationWithSpecifiedSource;
	---Purpose: Returns a ProductDefinitionFormationWithSpecifiedSource


	Init (me : mutable;
	      aId : mutable HAsciiString from TCollection;
	      aDescription : mutable HAsciiString from TCollection;
	      aOfProduct : mutable Product from StepBasic) is redefined;

	Init (me : mutable;
	      aId : mutable HAsciiString from TCollection;
	      aDescription : mutable HAsciiString from TCollection;
	      aOfProduct : mutable Product from StepBasic;
	      aMakeOrBuy : Source from StepBasic) is virtual;

	-- Specific Methods for Field Data Access --

	SetMakeOrBuy(me : mutable; aMakeOrBuy : Source);
	MakeOrBuy (me) returns Source;

fields

	makeOrBuy : Source from StepBasic; -- an Enumeration

end ProductDefinitionFormationWithSpecifiedSource;
