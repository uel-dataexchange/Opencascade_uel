-- File:	PColPGeom.cdl
-- Created:	Thu Jun  3 16:46:15 1993
-- Author:	fid
--		<model@mastox>
-- Copyright:	 Matra Datavision 1993


package PColPGeom 

        ---Purpose : This package  is used to  instantiate of  several
        --         generic classes from  the package  PCollection with
        --         objects from the package PGeom.

uses PCollection, PGeom

is


    class HArray1OfCurve 
    	instantiates HArray1 from PCollection (Curve from PGeom);
    class HArray1OfBoundedCurve 
    	instantiates HArray1 from PCollection (BoundedCurve from PGeom);
    class HArray1OfBezierCurve 
    	instantiates HArray1 from PCollection (BezierCurve from PGeom);
    class HArray1OfBSplineCurve 
    	instantiates HArray1 from PCollection (BSplineCurve from PGeom);
    class HArray1OfSurface 
    	instantiates HArray1 from PCollection (Surface from PGeom);
    class HArray1OfBoundedSurface 
    	instantiates HArray1 from PCollection (BoundedSurface from PGeom);



    class HArray2OfSurface 
    	instantiates HArray2 from PCollection (Surface from PGeom);
    class HArray2OfBoundedSurface 
    	instantiates HArray2 from PCollection (BoundedSurface from PGeom);
    class HArray2OfBezierSurface 
    	instantiates HArray2 from PCollection (BezierSurface from PGeom);
    class HArray2OfBSplineSurface 
    	instantiates HArray2 from PCollection (BSplineSurface from PGeom);



--    class HSequenceOfCurve  
--    	instantiates HSequence from PCollection (Curve from PGeom);
--    class HSequenceOfBoundedCurve  
--    	instantiates HSequence from PCollection (BoundedCurve from PGeom);
--    class HSequenceOfSurface 
--    	instantiates HSequence from PCollection (Surface from PGeom);
--    class HSequenceOfBoundedSurface 
--    	instantiates HSequence from PCollection (BoundedSurface from PGeom);


end PColPGeom;
