-- File:	RWStepBasic_RWMassUnit.cdl
-- Created:	Thu Dec 12 15:38:08 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWMassUnit from RWStepBasic

    ---Purpose: Read & Write tool for MassUnit

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    MassUnit from StepBasic

is
    Create returns RWMassUnit from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : MassUnit from StepBasic);
	---Purpose: Reads MassUnit

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: MassUnit from StepBasic);
	---Purpose: Writes MassUnit

    Share (me; ent : MassUnit from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWMassUnit;
