-- File:        PS_Driver.cdl
-- Created:     Tue Feb 22 08:46:41 1994
-- Author:      Jean Louis FRENKEL
--              <jlf@minox>
---Copyright:    Matra Datavision 1994

class Driver from PS inherits PlotterDriver from PlotMgt
  ---Purpose: This class defines a PS (Adobe PostScript) plotter Driver.
  ---         All necessary information about methods (purpose, level, category, etc.)
  ---         can be found in CDL files from the inheritance tree (PlotMgt_PlotterDriver,
  ---         Aspect_Driver).


uses
  Plotter            from PlotMgt,
  TypeOfColorSpace   from Aspect,
  FormatOfSheetPaper from Aspect,
  ExtendedString     from TCollection,
  AsciiString        from TCollection,
  ColorMap           from Aspect,
  TypeMap            from Aspect,
  WidthMap           from Aspect,
  FontMap            from Aspect,
  MarkMap            from Aspect,
  TypeOfText         from Aspect,
  TypeOfPrimitive    from Aspect,
  PlaneAngle         from Quantity,
  Length             from Quantity,
  Factor             from Quantity,
  Ratio              from Quantity


raises
  DriverError from Aspect


is
  Create(aName: CString from Standard;                   
      aDX,aDY: Length from Quantity;
      aTypeOfColorSpace: TypeOfColorSpace from Aspect = Aspect_TOCS_RGB;                 
      aSheetFormat: FormatOfSheetPaper from Aspect = Aspect_FOSP_A4)
  returns mutable Driver from PS;

  
  Create(aPlotter : Plotter from PlotMgt;
      aName: CString from Standard;       
      aPaperX,aPaperY: Length from Quantity;
      aTypeOfColorSpace: TypeOfColorSpace from Aspect = Aspect_TOCS_RGB)
  returns mutable Driver from PS;
---Purpose: Constructs a file called aName as the graphic
-- plotter file. The parameters of the plotter aPlotter
-- are taken into account for defining this plotter file.
-- aPaperX,aPaperY defines the size of the
-- sheet-paper and the value of aTypeOfColorSpace
-- defines the mode for processing colors.
  
  BeginFile(me: mutable;
          aPlotter : Plotter from PlotMgt;
          aName: CString from Standard;
          aDX,aDY: Length from Quantity;
          aTypeOfColorSpace: TypeOfColorSpace from Aspect;               
          aPaperX,aPaperY: Length from Quantity)
  is private;

  BeginDraw (me: mutable) is static;

---Purpose:
-- Begins a new page of graphics in the plotter file called "aName".
  EndDraw (me: mutable; dontFlush: Boolean = Standard_False) is static;


  ---------------------------------------------
  -- Category: Methods to define the attributes
  ---------------------------------------------
  InitializeColorMap(me: mutable; aColorMap: ColorMap from Aspect) 
  is virtual protected;


  InitializeTypeMap(me: mutable; aTypeMap: TypeMap from Aspect)
  is virtual protected;


  InitializeWidthMap(me: mutable; aWidthMap: WidthMap from Aspect)
  is virtual protected;


  InitializeFontMap(me: mutable; aFontMap: FontMap from Aspect)
  is virtual protected;


  InitializeMarkMap(me: mutable; aFontMap: MarkMap from Aspect)
  is virtual protected;


  ---------------------------------------------
  -- Category: Methods to set the attributes
  ---------------------------------------------
  SetTextAttrib (me: mutable;
     ColorIndex: Integer from Standard;
     FontIndex: Integer from Standard)
  is redefined;


  SetTextAttrib (me: mutable;
     ColorIndex: Integer from Standard;
     FontIndex: Integer from Standard;
     aSlant: PlaneAngle from Quantity;
     aHScale: Factor from Quantity;
     aWScale: Factor from Quantity;
     isUnderlined: Boolean from Standard = Standard_False)
  is redefined;


  --------------------------------
  -- Actual set graphic attributes
  --------------------------------
  PlotLineAttrib (me: mutable;
      ColorIndex: Integer from Standard;
      TypeIndex: Integer from Standard;
      WidthIndex: Integer from Standard)
  is redefined protected;


  -----------------------------------------
  -- Category: Methods to manage the images
  -----------------------------------------
  SizeOfImageFile (me; anImageFile: CString from Standard;
                       aWidth,aHeight: out Integer from Standard)
  returns Boolean from Standard is redefined;


  -----------------------------------------------
  -- Category: Private methods to draw primitives
  -----------------------------------------------
  PlotPoint (me : mutable; X, Y: ShortReal from Standard)
  returns Boolean from Standard
  is redefined protected;


  PlotSegment (me : mutable;
      X1, Y1: ShortReal from Standard;
      X2, Y2: ShortReal from Standard)
  returns Boolean from Standard
  is redefined protected;


  PlotPolyline (me : mutable;
      xArray : Address from Standard;
      yArray : Address from Standard;
      nPts   : Address from Standard;
      nParts : Integer from Standard)
  returns Boolean from Standard
  is redefined protected;


  PlotPolygon (me : mutable;
      xArray : Address from Standard;
      yArray : Address from Standard;
      nPts   : Address from Standard;
      nParts : Integer from Standard)
  returns Boolean from Standard
  is redefined protected;


  PlotArc (me : mutable; X,Y : ShortReal from Standard;
      anXradius,anYradius : ShortReal from Standard;
      sAngle: ShortReal from Standard;
      oAngle: ShortReal from Standard)
  returns Boolean from Standard
  is redefined protected;


  PlotPolyArc (me : mutable; X,Y : ShortReal from Standard;
      anXradius,anYradius : ShortReal from Standard;
      sAngle: ShortReal from Standard;
      oAngle: ShortReal from Standard)
  returns Boolean from Standard
  is redefined protected;


  PlotMarker (me : mutable;
      aMarker: Integer from Standard;
      Xpos:  ShortReal from Standard;
      Ypos:  ShortReal from Standard;
      Width: ShortReal from Standard;
      Height: ShortReal from Standard;
      Angle: ShortReal from Standard)
  returns Boolean from Standard
  is redefined protected;


  PlotText (me : mutable;
      aText: ExtendedString from TCollection;
      Xpos:  ShortReal from Standard;
      Ypos:  ShortReal from Standard;
      anAngle: ShortReal from Standard;
      aType: TypeOfText from Aspect)
  returns Boolean from Standard
  is redefined protected;
      

  PlotText (me : mutable;
      aText: CString from Standard;
      Xpos:  ShortReal from Standard;
      Ypos:  ShortReal from Standard;
      anAngle: ShortReal from Standard;
      aType: TypeOfText from Aspect)
  returns Boolean from Standard
  is redefined protected;


  PlotPolyText (me : mutable;
      aText: ExtendedString from TCollection;
      Xpos:  ShortReal from Standard;
      Ypos:  ShortReal from Standard;
      aMargin: Ratio from Quantity;
      anAngle: ShortReal from Standard;
      aType: TypeOfText from Aspect)
  returns Boolean from Standard
  is redefined protected;


  PlotPolyText (me : mutable;
      aText: CString from Standard;
      Xpos:  ShortReal from Standard;
      Ypos:  ShortReal from Standard;
      aMargin: Ratio from Quantity;
      anAngle: ShortReal from Standard;
      aType: TypeOfText from Aspect)
  returns Boolean from Standard
  is redefined protected;


  PlotImage (me: mutable; 
      aX, aY, aWidth:  ShortReal from Standard;
      aHeight, aScale: ShortReal from Standard;
      anImageFile:     CString   from Standard;
      anArrayOfPixels: Address   from Standard;
      aLineIndex:      Integer   from Standard = -1)
  returns Boolean from Standard
  is redefined protected;


  ----------------------------
  -- Category: Inquire methods
  ----------------------------
  Convert(me; aShortReal: ShortReal from Standard) 
  returns ShortReal from Standard is static private;
---Purpose: For this driver
-- - returns the DPU (device plotter unit) value
--   corresponding to the number of pixels PV, or
-- - returns the number of pixels corresponding to the DPU value DV, or
-- - returns the DPU coordinates (DX,DY)
--   corresponding to the pixel position (PX,PY), or
-- - returns the pixel position (PX,PY) corresponding to
--   the DPU coordinates (DX,DY).
--   The DPU value is specified in millimeters by default.
-- Warning
-- The pixel size is 325mm/1152 by default and can be
-- changed with the SetPixelSize function.

  DrawCurveCapable (me)
  returns Boolean from Standard is redefined protected;

  MapX(me; aShortReal: ShortReal from Standard) 
  returns ShortReal from Standard is redefined private;

  
  MapY(me; aShortReal: ShortReal from Standard) 
  returns ShortReal from Standard is redefined private; 

   
fields
  myCurrentPage: Integer from Standard;

end Driver from PS;
