-- File:	StepAP203_ContractedItem.cdl
-- Created:	Fri Nov 26 16:26:26 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class ContractedItem from StepAP203
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type ContractedItem

uses
    ProductDefinitionFormation from StepBasic

is
    Create returns ContractedItem from StepAP203;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of ContractedItem select type
	--          1 -> ProductDefinitionFormation from StepBasic
	--          0 else

    ProductDefinitionFormation (me) returns ProductDefinitionFormation from StepBasic;
	---Purpose: Returns Value as ProductDefinitionFormation (or Null if another type)

end ContractedItem;
