-- File:	IGESDimen_ToolDimensionedGeometry.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolDimensionedGeometry  from IGESDimen

    ---Purpose : Tool to work on a DimensionedGeometry. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses DimensionedGeometry from IGESDimen,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolDimensionedGeometry;
    ---Purpose : Returns a ToolDimensionedGeometry, ready to work


    ReadOwnParams (me; ent : mutable DimensionedGeometry;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : DimensionedGeometry;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : DimensionedGeometry;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a DimensionedGeometry <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable DimensionedGeometry) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a DimensionedGeometry
    --           (NbDimensions forced to 1)

    DirChecker (me; ent : DimensionedGeometry) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : DimensionedGeometry;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : DimensionedGeometry; entto : mutable DimensionedGeometry;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : DimensionedGeometry;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolDimensionedGeometry;
