-- File:        ReparametrisedCompositeCurveSegment.cdl
-- Created:     Fri Dec  1 11:11:26 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class ReparametrisedCompositeCurveSegment from StepGeom 

inherits CompositeCurveSegment from StepGeom 

uses

	Real from Standard, 
	TransitionCode from StepGeom, 
	Boolean from Standard, 
	Curve from StepGeom
is

	Create returns mutable ReparametrisedCompositeCurveSegment;
	---Purpose: Returns a ReparametrisedCompositeCurveSegment


	Init (me : mutable;
	      aTransition : TransitionCode from StepGeom;
	      aSameSense : Boolean from Standard;
	      aParentCurve : mutable Curve from StepGeom) is redefined;

	Init (me : mutable;
	      aTransition : TransitionCode from StepGeom;
	      aSameSense : Boolean from Standard;
	      aParentCurve : mutable Curve from StepGeom;
	      aParamLength : Real from Standard) is virtual;

	-- Specific Methods for Field Data Access --

	SetParamLength(me : mutable; aParamLength : Real);
	ParamLength (me) returns Real;

fields

	paramLength : Real from Standard;

end ReparametrisedCompositeCurveSegment;
