-- File:        DraughtingPreDefinedCurveFont.cdl
-- Created:     Mon Dec  4 12:02:25 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWDraughtingPreDefinedCurveFont from RWStepVisual

	---Purpose : Read & Write Module for DraughtingPreDefinedCurveFont

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     DraughtingPreDefinedCurveFont from StepVisual

is

	Create returns RWDraughtingPreDefinedCurveFont;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable DraughtingPreDefinedCurveFont from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : DraughtingPreDefinedCurveFont from StepVisual);

end RWDraughtingPreDefinedCurveFont;
