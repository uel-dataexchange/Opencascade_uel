-- File:	TopOpeBRepDS_FaceInterferenceTool.cdl
-- Created:	Tue Nov  8 14:47:14 1994
-- Author:	Jean Yves LEBEY
--		<jyl@bravox>
---Copyright:	 Matra Datavision 1994


class FaceInterferenceTool from TopOpeBRepDS 

---Purpose: a tool computing complex transition on Face.

uses

    Orientation from TopAbs,
    SurfaceTransition from TopTrans,
    Interference from TopOpeBRepDS,
    Curve from TopOpeBRepDS,
    Shape from TopoDS,
    Pnt from gp,
    Dir from gp,
    PDataStructure from TopOpeBRepDS
    
is

    Create(P : PDataStructure from TopOpeBRepDS)
    returns FaceInterferenceTool from TopOpeBRepDS;
    
    
    Init(me : in out; 
    	 FI : Shape from TopoDS; -- face accessing I
	 E : Shape from TopoDS; 
         Eisnew : Boolean;
         I : Interference from TopOpeBRepDS)
    ---Purpose: 
    -- Eisnew = true if E is a new edge built on edge I->Geometry()
    -- 	        false if E is shape <=> I->Geometry()
    is static;

    Add(me : in out;
    	FI : Shape from TopoDS; -- face accessing I
    	F : Shape from TopoDS;
	E : Shape from TopoDS;Eisnew : Boolean;
        I : Interference from TopOpeBRepDS)
    ---Purpose: 
    -- Eisnew = true if E is a new edge built on edge I->Geometry()
    -- 	        false if E is shape <=> I->Geometry()
    is static;
    
    Add(me : in out; 
        E : Shape from TopoDS;
	C : Curve from TopOpeBRepDS;
        I : Interference from TopOpeBRepDS)
    is static;

    SetEdgePntPar(me : in out; P : Pnt from gp; par : Real);
    GetEdgePntPar(me ; P : out Pnt from gp; par : out Real);
    IsEdgePntParDef(me) returns Boolean;

    Transition(me; I : mutable Interference from TopOpeBRepDS)
    is static;
    
fields
    
    myPBDS            : PDataStructure from TopOpeBRepDS; 
    myrefdef          : Boolean; -- myTool has been initialized   
    myFaceOrientation : Orientation from TopAbs;
    myFaceOriented    : Integer from Standard;
    myTool            : SurfaceTransition from TopTrans;
    myEdge            : Shape from TopoDS;  -- geometric domain where happens the interference
    isLine            : Boolean;
    myPntOnEd         : Pnt from gp; -- point on edge where is locally described the interference.
    myParOnEd         : Real;        -- point parameter on edge.
    myOnEdDef         : Boolean;
    myTole            : Real; 


end FaceInterferenceTool from TopOpeBRepDS;
