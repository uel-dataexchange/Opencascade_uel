-- File:	StepFEA_CurveElementIntervalLinearlyVarying.cdl
-- Created:	Wed Jan 22 17:31:43 2003 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class CurveElementIntervalLinearlyVarying from StepFEA
inherits CurveElementInterval from StepFEA

    ---Purpose: Representation of STEP entity CurveElementIntervalLinearlyVarying

uses
    CurveElementLocation from StepFEA,
    EulerAngles from StepBasic,
    HArray1OfCurveElementSectionDefinition from StepElement

is
    Create returns CurveElementIntervalLinearlyVarying from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aCurveElementInterval_FinishPosition: CurveElementLocation from StepFEA;
                       aCurveElementInterval_EuAngles: EulerAngles from StepBasic;
                       aSections: HArray1OfCurveElementSectionDefinition from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    Sections (me) returns HArray1OfCurveElementSectionDefinition from StepElement;
	---Purpose: Returns field Sections
    SetSections (me: mutable; Sections: HArray1OfCurveElementSectionDefinition from StepElement);
	---Purpose: Set field Sections

fields
    theSections: HArray1OfCurveElementSectionDefinition from StepElement;

end CurveElementIntervalLinearlyVarying;
