-- File:	MDataXtd_PatternStdRetrievalDriver.cdl
-- Created:	Mon Feb 16 14:33:53 1998
-- Author:	Jing Cheng MEI
--		<mei@pinochiox.paris1.matra-dtv.fr>
-- modified     Sergey Zaritchny
---Copyright:	 Matra Datavision 1998

class PatternStdRetrievalDriver from MDataXtd  inherits ARDriver from MDF

	---Purpose: 

uses RRelocationTable from MDF,
     Attribute        from PDF,
     Attribute        from TDF, 
     MessageDriver    from CDM

is


    Create(theMessageDriver : MessageDriver from CDM)  -- Version 0
    returns mutable PatternStdRetrievalDriver from MDataXtd;
    

    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type: PatternStd from PDataXtd.

    NewEmpty (me)  returns mutable Attribute from TDF;


    Paste(me;
    	  Source     :         Attribute from PDF;
    	  Target     : mutable Attribute from TDF;
    	  RelocTable : RRelocationTable  from MDF);

end PatternStdRetrievalDriver;

