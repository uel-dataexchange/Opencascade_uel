-- File:	StepBasic_GroupRelationship.cdl
-- Created:	Wed May 10 15:09:07 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class GroupRelationship from StepBasic
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity GroupRelationship

uses
    HAsciiString from TCollection,
    Group from StepBasic

is
    Create returns GroupRelationship from StepBasic;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       hasDescription: Boolean;
                       aDescription: HAsciiString from TCollection;
                       aRelatingGroup: Group from StepBasic;
                       aRelatedGroup: Group from StepBasic);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description
    HasDescription (me) returns Boolean;
	---Purpose: Returns True if optional field Description is defined

    RelatingGroup (me) returns Group from StepBasic;
	---Purpose: Returns field RelatingGroup
    SetRelatingGroup (me: mutable; RelatingGroup: Group from StepBasic);
	---Purpose: Set field RelatingGroup

    RelatedGroup (me) returns Group from StepBasic;
	---Purpose: Returns field RelatedGroup
    SetRelatedGroup (me: mutable; RelatedGroup: Group from StepBasic);
	---Purpose: Set field RelatedGroup

fields
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection; -- optional
    theRelatingGroup: Group from StepBasic;
    theRelatedGroup: Group from StepBasic;
    defDescription: Boolean; -- flag "is Description defined"

end GroupRelationship;
