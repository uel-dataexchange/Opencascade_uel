-- File:	Graphic3d_ArrayOfQuadrangles.cdl
-- Created:	04/01/01 : GG : G005 : Draw ARRAY primitives
--

class ArrayOfQuadrangles from Graphic3d inherits ArrayOfPrimitives from Graphic3d 

uses
	Color			from Quantity,
	Pnt			from gp,
	Pnt2d			from gp,
	Dir			from gp

raises
    OutOfRange from Standard

is

	-- constructor
	Create (
                maxVertexs: Integer from Standard;
                maxEdges: Integer from Standard = 0;
                hasVNormals: Boolean from Standard = Standard_False;
                hasVColors: Boolean from Standard = Standard_False;
                hasTexels: Boolean from Standard = Standard_False;
		hasEdgeInfos: Boolean from Standard = Standard_False)
	returns mutable ArrayOfQuadrangles from Graphic3d;
        ---Purpose: Creates an array of quadrangles,
	-- a quadrangle can be filled as:
	-- 1) creating a set of quadrangles defined with his vertexs.
	--    i.e:
	--    myArray = Graphic3d_ArrayOfQuadrangles(8)
	--    myArray->AddVertex(x1,y1,z1) 
	--	....
	--    myArray->AddVertex(x8,y8,z8) 
	-- 3) creating a set of indexed quadrangles defined with his vertex
	--    ans edges. 
	--    i.e:
	--    myArray = Graphic3d_ArrayOfQuadrangles(6,8)
	--    myArray->AddVertex(x1,y1,z1) 
	--	....
	--    myArray->AddVertex(x6,y6,z6) 
	--    myArray->AddEdge(1)
	--    myArray->AddEdge(2)
	--    myArray->AddEdge(3)
	--    myArray->AddEdge(4)
	--    myArray->AddEdge(3)
	--    myArray->AddEdge(4)
	--    myArray->AddEdge(5)
	--    myArray->AddEdge(6)
	-- 
	-- <maxVertexs> defined the maximun allowed vertex number in the array.
	-- <maxEdges> defined the maximun allowed edge number in the array.
	--  Warning:
	-- When <hasVNormals> is TRUE , you must use one of
	--	AddVertex(Point,Normal) 
	--  or  AddVertex(Point,Normal,Color)
	--  or  AddVertex(Point,Normal,Texel) methods.
	-- When <hasVColors> is TRUE , you must use one of
	--	AddVertex(Point,Color)
	--  or  AddVertex(Point,Normal,Color) methods.
	-- When <hasTexels> is TRUE , you must use one of
	--	AddVertex(Point,Texel) 
	--  or  AddVertex(Point,Normal,Texel) methods.
	-- When <hasEdgeInfos> is TRUE , <maxEdges> must be > 0 and
	--	you must use the
	--	AddEdge(number,visibillity) method.
	--  Warning:
	-- the user is responsible about the orientation of the quadrangle
	-- depending of the order of the created vertex or edges and this
	-- orientation must be coherent with the vertex normal optionnaly
	-- given at each vertex (See the Orientate() methods).

end;
