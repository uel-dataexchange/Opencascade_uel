-- File:	Voxel_OctBoolDS.cdl
-- Created:	Sun Aug 26 12:21:23 2008
-- Author:	Vladislav ROMASHKO
--		<vladislav.romashko@opencascade.com>
---Copyright:	Open CASCADE S.A.

class OctBoolDS from Voxel inherits DS from Voxel

    ---Purpose: A 3D voxel model keeping a boolean flag (1 or 0)
    --          value for each voxel, and having an opportunity to split each voxel
    --          into 8 sub-voxels.

is

    Create
    ---Purpose: An empty constructor.
    returns OctBoolDS from Voxel;

    Create(x     : Real    from Standard;
    	   y     : Real    from Standard;
    	   z     : Real    from Standard;
    	   x_len : Real    from Standard;
    	   y_len : Real    from Standard;
    	   z_len : Real    from Standard;
	   nb_x  : Integer from Standard;
	   nb_y  : Integer from Standard;
	   nb_z  : Integer from Standard)
    ---Purpose: A constructor initializing the voxel model.
    --          (x, y, z) - the start point of the box.
    --          (x_len, y_len, z_len) - lengths in x, y and z directions along axes of a co-ordinate system.
    --          (nb_x, nb_y, nb_z) - number of splits (voxels) along x, y and z directions.
    returns OctBoolDS from Voxel;

    Init(me : in out;
    	 x     : Real    from Standard;
    	 y     : Real    from Standard;
    	 z     : Real    from Standard;
    	 x_len : Real    from Standard;
    	 y_len : Real    from Standard;
    	 z_len : Real    from Standard;
	 nb_x  : Integer from Standard;
	 nb_y  : Integer from Standard;
	 nb_z  : Integer from Standard)
    ---Purpose: Initialization of the voxel model.
    --          (x, y, z) - the start point of the box.
    --          (x_len, y_len, z_len) - lengths in x, y and z directions along axes of a co-ordinate system.
    --          (nb_x, nb_y, nb_z) - number of splits (voxels) along x, y and z directions.
    is redefined virtual;

    Destroy(me : in out);
    ---C++: alias ~
    ---Purpose: A destructor of the voxel model.

    SetZero(me : in out);
    ---Purpose: The method sets all values equal to 0 (false) and
    --          releases the memory.

    OptimizeMemory(me : in out);
    ---Purpose: The method searches voxels with equal-value of sub-voxels
    --          and removes them (remaining the value for the voxel).

    Set(me   : in out;
    	ix   : Integer from Standard;
    	iy   : Integer from Standard;
    	iz   : Integer from Standard;
	data : Boolean from Standard);
    ---Purpose: Defines a value for voxel with co-ordinates (ix, iy, iz).
    --          If the voxel is split into 8 sub-voxels, the split disappears.
    --          Initial state of the model is so that all voxels have value 0 (false),
    --          and this data doesn't occupy memory.
    --          Memory for data is allocating during setting non-zero values (true).

    Set(me   : in out;
    	ix   : Integer from Standard;
    	iy   : Integer from Standard;
    	iz   : Integer from Standard;
	ioct : Integer from Standard;
	data : Boolean from Standard);
    ---Purpose: Defines a value for a sub-voxel of a voxel with co-ordinates (ix, iy, iz).
    --          If the voxel is not split into 8 sub-voxels yet, this method splits the voxel.
    --          Range of sub-voxels is 0 - 7.

    Get(me;
    	ix : Integer from Standard;
    	iy : Integer from Standard;
    	iz : Integer from Standard)
    ---Purpose: Returns the value of voxel with co-ordinates (ix, iy, iz).
    --          Warning!: the returned value may not coincide with the value of its 8 sub-voxels.
    --          Use the method ::IsSplit() to check whether a voxel has sub-voxels.
    returns Boolean from Standard;

    Get(me;
    	ix   : Integer from Standard;
    	iy   : Integer from Standard;
    	iz   : Integer from Standard;
    	ioct : Integer from Standard)
    ---Purpose: Returns the value of a sub-voxel of a voxel with co-ordinates (ix, iy, iz).
    --          If the voxel is not split, it returns the value of the voxel.
    --          Range of sub-voxels is 0 - 7.
    returns Boolean from Standard;

    IsSplit(me;
    	    ix   : Integer from Standard;
    	    iy   : Integer from Standard;
    	    iz   : Integer from Standard)
    ---Purpose: Returns true if the voxel is split into 8 sub-voxels.
    returns Boolean from Standard;


    ---Category: Private area
    --           ============

    Split(me : in out;
    	  ix   : Integer from Standard;
    	  iy   : Integer from Standard;
    	  iz   : Integer from Standard)
    is private;

    UnSplit(me : in out;
    	    ix   : Integer from Standard;
    	    iy   : Integer from Standard;
    	    iz   : Integer from Standard)
    is private;


fields

    mySubVoxels : Address from Standard;

end OctBoolDS;
