-- File:	RWStepRepr_RWShapeAspectRelationship.cdl
-- Created:	Tue Apr 18 16:42:58 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWShapeAspectRelationship from RWStepRepr

    ---Purpose: Read & Write tool for ShapeAspectRelationship

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ShapeAspectRelationship from StepRepr

is
    Create returns RWShapeAspectRelationship from RWStepRepr;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ShapeAspectRelationship from StepRepr);
	---Purpose: Reads ShapeAspectRelationship

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ShapeAspectRelationship from StepRepr);
	---Purpose: Writes ShapeAspectRelationship

    Share (me; ent : ShapeAspectRelationship from StepRepr;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWShapeAspectRelationship;
