-- File:	StepElement_ElementDescriptor.cdl
-- Created:	Thu Dec 12 17:29:00 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class ElementDescriptor from StepElement
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity ElementDescriptor

uses
    ElementOrder from StepElement,
    HAsciiString from TCollection

is
    Create returns ElementDescriptor from StepElement;
	---Purpose: Empty constructor

    Init (me: mutable; aTopologyOrder: ElementOrder from StepElement;
                       aDescription: HAsciiString from TCollection);
	---Purpose: Initialize all fields (own and inherited)

    TopologyOrder (me) returns ElementOrder from StepElement;
	---Purpose: Returns field TopologyOrder
    SetTopologyOrder (me: mutable; TopologyOrder: ElementOrder from StepElement);
	---Purpose: Set field TopologyOrder

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description

fields
    theTopologyOrder: ElementOrder from StepElement;
    theDescription: HAsciiString from TCollection;

end ElementDescriptor;
