-- File:	RWStepElement_RWSurfaceSectionField.cdl
-- Created:	Thu Dec 12 17:29:04 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWSurfaceSectionField from RWStepElement

    ---Purpose: Read & Write tool for SurfaceSectionField

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    SurfaceSectionField from StepElement

is
    Create returns RWSurfaceSectionField from RWStepElement;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : SurfaceSectionField from StepElement);
	---Purpose: Reads SurfaceSectionField

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: SurfaceSectionField from StepElement);
	---Purpose: Writes SurfaceSectionField

    Share (me; ent : SurfaceSectionField from StepElement;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWSurfaceSectionField;
