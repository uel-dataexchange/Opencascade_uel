-- File:	GeomToStep_MakeSurface.cdl
-- Created:	Tue Jun 22 12:19:43 1993
-- Author:	Martine LANGLOIS
--		<mla@mastox>
---Copyright:	 Matra Datavision 1993

class MakeSurface from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          Surface from Geom and the class Surface from StepGeom which
    --          describes a Surface from prostep. As Surface is an abstract
    --          Surface this class is an access to the sub-class required.
  
uses Surface from Geom,
     Surface from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( C : Surface from Geom ) returns MakeSurface;

Value (me) returns Surface from StepGeom
    raises NotDone
    is static;
    ---C++: return const&

fields

    theSurface : Surface from StepGeom;
    	-- The solution from StepGeom
    	
end MakeSurface;



