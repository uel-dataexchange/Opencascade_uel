-- File:	StepFEA_ConstantSurface3dElementCoordinateSystem.cdl
-- Created:	Thu Dec 26 15:06:35 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class ConstantSurface3dElementCoordinateSystem from StepFEA
inherits FeaRepresentationItem from StepFEA

    ---Purpose: Representation of STEP entity ConstantSurface3dElementCoordinateSystem

uses
    HAsciiString from TCollection

is
    Create returns ConstantSurface3dElementCoordinateSystem from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aAxis: Integer;
                       aAngle: Real);
	---Purpose: Initialize all fields (own and inherited)

    Axis (me) returns Integer;
	---Purpose: Returns field Axis
    SetAxis (me: mutable; Axis: Integer);
	---Purpose: Set field Axis

    Angle (me) returns Real;
	---Purpose: Returns field Angle
    SetAngle (me: mutable; Angle: Real);
	---Purpose: Set field Angle

fields
    theAxis: Integer;
    theAngle: Real;

end ConstantSurface3dElementCoordinateSystem;
