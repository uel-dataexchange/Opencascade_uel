-- File:	Quantity_Convert.cdl
-- Created:	Tue Jul 19 16:36:20 1994
-- Author:	Guest Kernel
--		<g_kernel@bibox>
---Copyright:	 Matra Datavision 1994


class Convert from Quantity

    	---Purpose: Services to manage units conversion between Front-ends and Engines.
    	-- This conversion is managed by a table of correspondance between the quantities
    	-- and their "conversion coefficient".
    	-- This table is implemented like an external array (TCollection_Array1) regarding 
    	-- to the quantities enumeration.
     
uses 
    AsciiString from TCollection,
    PhysicalQuantity from Quantity,
    Coefficient from Quantity
	     
is

    Create returns Convert from Quantity;
    	---Purpose: Creates an object;

    SetQuantity(myclass ; 
                aQuantity : PhysicalQuantity from Quantity ;
	        aCoef: Coefficient from Quantity);	    
    	---Purpose: Updates the conversion table (correspondances between 
    	-- Quantities and conversion coefficients).
    	---C++: inline

    ConvertUserToSI(myclass ; 
                    aQuantity : PhysicalQuantity from Quantity ;
          	    aVal : Real from Standard)
    returns Real from Standard;
        ---Purpose: Converts, from the conversion table, the value <aVal>
    	-- from the user system to the SI system. 
    	---C++: inline

    ConvertSIToUser(myclass ; 
                    aQuantity : PhysicalQuantity from Quantity ;
          	    aVal : Real from Standard)
    returns Real from Standard;
    	---Purpose: Converts, from the conversion table, the value <aVal>
   	-- from the SI system to the user system. 
    	---C++: inline

    IsPhysicalQuantity(myclass; 
                       aTypeName : AsciiString from TCollection ; 
                       anEnum : in out AsciiString from TCollection)
    returns Boolean from Standard;
    	---Purpose:
    	-- if (aType is a physical quantity)
    	--    returns True and the name of the associated PhysicalQuantity .
    	-- else 
    	--    returns False.

end Convert from Quantity;
	        	







































































































