-- File:	IGESDefs_ToolGenericData.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolGenericData  from IGESDefs

    ---Purpose : Tool to work on a GenericData. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses GenericData from IGESDefs,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolGenericData;
    ---Purpose : Returns a ToolGenericData, ready to work


    ReadOwnParams (me; ent : mutable GenericData;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : GenericData;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : GenericData;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a GenericData <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : GenericData) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : GenericData;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : GenericData; entto : mutable GenericData;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : GenericData;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolGenericData;
