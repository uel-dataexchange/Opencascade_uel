-- File:	RWStepBasic_RWObjectRole.cdl
-- Created:	Wed May 10 15:09:08 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWObjectRole from RWStepBasic

    ---Purpose: Read & Write tool for ObjectRole

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ObjectRole from StepBasic

is
    Create returns RWObjectRole from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ObjectRole from StepBasic);
	---Purpose: Reads ObjectRole

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ObjectRole from StepBasic);
	---Purpose: Writes ObjectRole

    Share (me; ent : ObjectRole from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWObjectRole;
