-- File:        OrganizationalAddress.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWOrganizationalAddress from RWStepBasic

	---Purpose : Read & Write Module for OrganizationalAddress

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     OrganizationalAddress from StepBasic,
     EntityIterator from Interface

is

	Create returns RWOrganizationalAddress;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable OrganizationalAddress from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : OrganizationalAddress from StepBasic);

	Share(me; ent : OrganizationalAddress from StepBasic; iter : in out EntityIterator);

end RWOrganizationalAddress;
