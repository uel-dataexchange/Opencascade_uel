-- File:	IGESSelect_UpdateLastChange.cdl
-- Created:	Wed Jun  1 16:19:53 1994
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1994


class UpdateLastChange  from IGESSelect  inherits ModelModifier from IGESSelect

    ---Purpose : Allows to Change the Last Change Date indication in the Header
    --           (Global Section) of IGES File. It is taken from the operating
    --           system (time of application of the Modifier).
    --           The Selection of the Modifier is not used : it simply acts as
    --           a criterium to select IGES Files to touch up.
    --           Remark : IGES Models noted as version before IGES 5.1 are in
    --           addition changed to 5.1

uses AsciiString from TCollection,
     IGESModel, CopyTool, ContextModif

is

    Create returns mutable UpdateLastChange;
    ---Purpose : Creates an UpdateLastChange, which uses the system Date

    Performing (me; ctx : in out ContextModif;
    	        target  : mutable IGESModel;
                TC      : in out CopyTool);
    ---Purpose : Specific action : only <target> is used : the system Date
    --           is set to Global Section Item n0 25. Also sets IGES Version
    --           (Item n0 23) to IGES5 if it was older.

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text which is
    --           "Update IGES Header Last Change Date"

end UpdateLastChange;
