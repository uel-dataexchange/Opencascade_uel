-- File:	MakeArcOfParabola.cdl
-- Created:	Mon Sep 28 11:51:03 1992
-- Author:	Remi GILET
--		<reg@sdsun2>
---Copyright:	 Matra Datavision 1992

class MakeArcOfParabola from GC inherits Root from GC
    	---Purpose: Implements construction algorithms for an arc
    	-- of parabola in 3D space. The result is a Geom_TrimmedCurve curve.
    	-- A MakeArcOfParabola object provides a framework for:
    	-- -   defining the construction of the arc of parabola,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the results. In particular, the
    	--   Value function returns the constructed arc of parabola.
uses Pnt          from gp,
     Parab        from gp,
     Dir          from gp,
     Ax1          from gp,
     Real         from Standard,
     TrimmedCurve from Geom

raises NotDone from StdFail

is

Create(Parab          : Parab   from gp       ;
       Alpha1, Alpha2 : Real    from Standard ;
       Sense          : Boolean from Standard ) returns MakeArcOfParabola;
    	---Purpose: Creates an arc of Parabola (TrimmedCurve from Geom) from 
    	--          a Parabola between two parameters Alpha1 and Alpha2
    	--          (given in radians).

Create(Parab : Parab   from gp       ;
       P     : Pnt     from gp       ;
       Alpha : Real    from Standard ;
       Sense : Boolean from Standard ) returns MakeArcOfParabola;
    	---Purpose: Creates an arc of Parabola (TrimmedCurve from Geom) from 
    	--          a Parabola between point <P> and the parameter
        --          Alpha (given in radians).

Create(Parab : Parab   from gp ;
       P1    : Pnt     from gp ;
       P2    : Pnt     from gp ;
       Sense : Boolean from Standard ) returns MakeArcOfParabola;
    	---Purpose: Creates an arc of Parabola (TrimmedCurve from Geom) from 
    	--          a Parabola between two points P1 and P2.

Value(me) returns TrimmedCurve from Geom
    raises NotDone
    is static;
    	---Purpose: Returns the constructed arc of parabola.
    	---C++: return const&

Operator(me) returns TrimmedCurve from Geom
    is static;
    	---C++: return const&
    	---C++: alias "Standard_EXPORT operator Handle_Geom_TrimmedCurve() const;"

fields

    TheArc : TrimmedCurve from Geom;
    --The solution from Geom.
    
end MakeArcOfParabola;
