-- File:	GraphTools_VertexIterator.cdl
-- Created:	Wed Mar  6 18:20:11 1991
-- Author:	Denis Pascal
--		<dp@topsn3>
---Copyright:	 Matra Datavision 1991, 1992


generic class VertexIterator from GraphTools (Graph  as any;
		    		               Vertex as any)
				  
--template class VertexIterator from GraphTools (Graph  as any,
--                                                 Vertex as any)
				  
    ---Purpose: Template class which  defines Signature of an iterator
    --          to visit each adjacent vertex  of a  given one  in the
    --          underlying graph.


raises NoMoreObject from Standard,
       NoSuchObject from Standard

is

    Create (G : Graph; V : Vertex) returns VertexIterator;

    More (me) returns Boolean;
	---Purpose: Returns TRUE if there are other vertices.
       ---Level: Public

    Next(me : in out)
    	--- Purpose : Set the iterator to the next Vertex.
       ---Level: Public
    raises NoMoreObject from Standard;

    Value(me) returns Vertex
	--- Purpose: Returns the vertex value for the current position
	--           of the iterator.
       ---Level: Public
    raises NoSuchObject from Standard;

end VertexIterator;



















