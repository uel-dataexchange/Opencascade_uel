-- File:	RWStepDimTol_RWCircularRunoutTolerance.cdl
-- Created:	Wed Jun  4 13:34:34 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWCircularRunoutTolerance from RWStepDimTol

    ---Purpose: Read & Write tool for CircularRunoutTolerance

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    CircularRunoutTolerance from StepDimTol

is
    Create returns RWCircularRunoutTolerance from RWStepDimTol;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : CircularRunoutTolerance from StepDimTol);
	---Purpose: Reads CircularRunoutTolerance

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: CircularRunoutTolerance from StepDimTol);
	---Purpose: Writes CircularRunoutTolerance

    Share (me; ent : CircularRunoutTolerance from StepDimTol;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWCircularRunoutTolerance;
