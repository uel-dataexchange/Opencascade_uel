-- File:	StepRepr_PropertyDefinition.cdl
-- Created:	Mon Jul  3 16:29:03 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class PropertyDefinition from StepRepr
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity PropertyDefinition

uses
    HAsciiString from TCollection,
    CharacterizedDefinition from StepRepr

is
    Create returns PropertyDefinition from StepRepr;
	---Purpose: Empty constructor

    Init (me: mutable; aName: HAsciiString from TCollection;
                       hasDescription: Boolean;
                       aDescription: HAsciiString from TCollection;
                       aDefinition: CharacterizedDefinition from StepRepr);
	---Purpose: Initialize all fields (own and inherited)

    Name (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Name
    SetName (me: mutable; Name: HAsciiString from TCollection);
	---Purpose: Set field Name

    Description (me) returns HAsciiString from TCollection;
	---Purpose: Returns field Description
    SetDescription (me: mutable; Description: HAsciiString from TCollection);
	---Purpose: Set field Description
    HasDescription (me) returns Boolean;
	---Purpose: Returns True if optional field Description is defined

    Definition (me) returns CharacterizedDefinition from StepRepr;
	---Purpose: Returns field Definition
    SetDefinition (me: mutable; Definition: CharacterizedDefinition from StepRepr);
	---Purpose: Set field Definition

fields
    theName: HAsciiString from TCollection;
    theDescription: HAsciiString from TCollection; -- optional
    theDefinition: CharacterizedDefinition from StepRepr;
    defDescription: Boolean; -- flag "is Description defined"

end PropertyDefinition;
