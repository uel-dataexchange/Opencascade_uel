-- File:        XmlMDataStd_VariableDriver.cdl
-- Created:     Fri Aug 24 20:16:51 2001
-- Author:      Alexander GRIGORIEV
-- Copyright:   Open Cascade 2001

class VariableDriver from XmlMDataStd  inherits ADriver from XmlMDF

        ---Purpose: Attribute Driver.

uses
    SRelocationTable from XmlObjMgt,
    RRelocationTable from XmlObjMgt,
    Persistent       from XmlObjMgt,
    MessageDriver    from CDM,
    Attribute        from TDF

is
    Create (theMessageDriver:MessageDriver from CDM)
        returns mutable VariableDriver from XmlMDataStd;

    NewEmpty (me)  returns mutable Attribute from TDF;

    Paste(me; Source     : Persistent from XmlObjMgt;
              Target     : mutable Attribute from TDF;
              RelocTable : out RRelocationTable from XmlObjMgt)
        returns Boolean from Standard;

    Paste(me; Source     : Attribute from TDF;
              Target     : in out Persistent from XmlObjMgt;
              RelocTable : out SRelocationTable from XmlObjMgt);

end VariableDriver;
