-- File:	RWStepBasic_RWIdentificationAssignment.cdl
-- Created:	Wed May 10 15:09:08 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWIdentificationAssignment from RWStepBasic

    ---Purpose: Read & Write tool for IdentificationAssignment

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    IdentificationAssignment from StepBasic

is
    Create returns RWIdentificationAssignment from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : IdentificationAssignment from StepBasic);
	---Purpose: Reads IdentificationAssignment

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: IdentificationAssignment from StepBasic);
	---Purpose: Writes IdentificationAssignment

    Share (me; ent : IdentificationAssignment from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWIdentificationAssignment;
