-- File:	Interface_Category.cdl
-- Created:	Wed Nov  8 19:11:08 1995
-- Author:	Christian CAILLET
--		<cky@fidox>
---Copyright:	 Matra Datavision 1995


class Category  from Interface

    ---Purpose : This class manages categories
    --           A category is defined by a name and a number, and can be
    --           seen as a way of rough classification, i.e. less precise than
    --           a cdl type.
    --           Hence, it is possible to dispatch every entity in about
    --           a dozen of categories, twenty is a reasonable maximum.
    --           
    --           Basically, the system provides the following categories :
    --           Shape (Geometry, BRep, CSG, Features, etc...)
    --           Drawing (Drawing, Views, Annotations, Pictures, Scketches ...)
    --           Structure (Component & Part, Groups & Patterns ...)
    --           Description (Meta-Data : Relations, Properties, Product ...)
    --           Auxiliary   (those which do not enter in the above list)
    --             and some dedicated categories
    --           FEA , Kinematics , Piping , etc...
    --           plus Professional  for other dedicated non-classed categories
    --           
    --           In addition, this class provides a way to compute then quickly
    --           query category numbers for an entire model.
    --           Values are just recorded as a list of numbers, control must
    --           then be done in a wider context (which must provide a Graph)

uses Integer, CString, Transient, HArray1OfInteger from TColStd,
     Protocol, GTool, InterfaceModel, ShareTool

is

    Create returns Category;
    ---Purpose : Creates a Category, with no protocol yet

    Create (proto : Protocol) returns Category;
    ---Purpose : Creates a Category with a given protocol

    Create (gtool : GTool) returns Category;
    ---Purpose : Creates a Category with a given GTool

    SetProtocol (me : in out; proto : Protocol);
    ---Purpose : Sets/Changes Protocol

    CatNum (me : in out; ent : Transient; shares : ShareTool)  returns Integer;
    ---Purpose : Determines the Category Number for an entity in its context,
    --           by using general service CategoryNumber

    ClearNums (me : in out);
    ---Purpose : Clears the recorded list of category numbers for a Model

    Compute  (me : in out; model : InterfaceModel; shares : ShareTool);
    ---Purpose : Computes the Category Number for each entity and records it,
    --           in an array (ent.number -> category number)
    --           Hence, it can be queried by the method Num.
    --           The Model itself is not recorded, this method is intended to
    --           be used in a wider context (which detains also a Graph, etc)

    Num (me; nument : Integer) returns Integer;
    ---Purpose : Returns the category number recorded for an entity number
    --           Returns 0 if out of range

    AddCategory (myclass; name : CString)  returns Integer;
    ---Purpose : Records a new Category defined by its names, produces a number
    --           New if not yet recorded

    NbCategories (myclass) returns Integer;
    ---Purpose : Returns the count of recorded categories

    Name (myclass; num : Integer) returns CString;
    ---Purpose : Returns the name of a category, according to its number

    Number (myclass; name : CString) returns Integer;
    ---Purpose : Returns the number of a category, according to its name


    Init (myclass);
    ---Purpose : Default initialisation
    --           (protected against several calls : passes only once)

fields

    thegtool : GTool;
    thenum   : HArray1OfInteger;

end Category;
