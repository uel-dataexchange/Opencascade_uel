-- File:        CompositeCurve.cdl
-- Created:     Fri Dec  1 11:11:16 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class CompositeCurve from StepGeom 

inherits BoundedCurve from StepGeom 

uses

	HArray1OfCompositeCurveSegment from StepGeom, 
	Logical from StepData, 
	CompositeCurveSegment from StepGeom, 
	HAsciiString from TCollection
is

	Create returns mutable CompositeCurve;
	---Purpose: Returns a CompositeCurve


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aSegments : mutable HArray1OfCompositeCurveSegment from StepGeom;
	      aSelfIntersect : Logical from StepData) is virtual;

	-- Specific Methods for Field Data Access --

	SetSegments(me : mutable; aSegments : mutable HArray1OfCompositeCurveSegment);
	Segments (me) returns mutable HArray1OfCompositeCurveSegment;
	SegmentsValue (me; num : Integer) returns mutable CompositeCurveSegment;
	NbSegments (me) returns Integer;
	SetSelfIntersect(me : mutable; aSelfIntersect : Logical);
	SelfIntersect (me) returns Logical;

fields

	segments : HArray1OfCompositeCurveSegment from StepGeom;
	selfIntersect : Logical from StepData;

end CompositeCurve;
