-- File:	RWStepBasic_RWDocument.cdl
-- Created:	Thu May 11 16:38:00 2000 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWDocument from RWStepBasic

    ---Purpose: Read & Write tool for Document

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    Document from StepBasic

is
    Create returns RWDocument from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : Document from StepBasic);
	---Purpose: Reads Document

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: Document from StepBasic);
	---Purpose: Writes Document

    Share (me; ent : Document from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWDocument;
