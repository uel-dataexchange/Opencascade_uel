-- File:	RWStepBasic_RWEffectivityAssignment.cdl
-- Created:	Wed May 10 15:09:06 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWEffectivityAssignment from RWStepBasic

    ---Purpose: Read & Write tool for EffectivityAssignment

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    EffectivityAssignment from StepBasic

is
    Create returns RWEffectivityAssignment from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : EffectivityAssignment from StepBasic);
	---Purpose: Reads EffectivityAssignment

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: EffectivityAssignment from StepBasic);
	---Purpose: Writes EffectivityAssignment

    Share (me; ent : EffectivityAssignment from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWEffectivityAssignment;
