-- File:	PTopoDS_Edge.cdl
-- Created:	Wed May  5 16:55:27 1993
-- Author:	Remi LEQUETTE
--		<rle@sdsun1>
---Copyright:	 Matra Datavision 1993



class Edge from PTopoDS inherits HShape from PTopoDS

is
    Create returns mutable Edge from PTopoDS;
	---Level: Internal 

end Edge;
