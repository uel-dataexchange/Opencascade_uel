-- File:	TPrsStd_NamedShapeDriver.cdl
-- Created:	Fri Aug  1 11:21:30 1997
-- Author:	SMO
---Copyright:	 Matra Datavision 1997


class NamedShapeDriver from TPrsStd inherits Driver from TPrsStd
---Purpose: An implementation of TPrsStd_Driver for named shapes.
uses

  GUID               from Standard,
  Label              from TDF,
  InteractiveObject  from AIS
is

    Create
    returns mutable NamedShapeDriver from TPrsStd;
---Purpose: Constructs an empty named shape driver.
    Update (me : mutable ;
           aLabel      : Label from TDF;
	   anAISObject : in out InteractiveObject from AIS)
    returns Boolean from Standard
    is  redefined virtual;
    --- Purpose: Build the AISObject (if null) or update it.
    --           No compute is done.
    --           Returns <True> if informations was found
    --           and AISObject updated. 
	   

end NamedShapeDriver;

