-- File:	RWStepFEA_RWFeaRepresentationItem.cdl
-- Created:	Thu Dec 12 17:51:06 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFeaRepresentationItem from RWStepFEA

    ---Purpose: Read & Write tool for FeaRepresentationItem

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FeaRepresentationItem from StepFEA

is
    Create returns RWFeaRepresentationItem from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FeaRepresentationItem from StepFEA);
	---Purpose: Reads FeaRepresentationItem

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FeaRepresentationItem from StepFEA);
	---Purpose: Writes FeaRepresentationItem

    Share (me; ent : FeaRepresentationItem from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFeaRepresentationItem;
