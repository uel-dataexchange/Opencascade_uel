-- File:	IGESSelect_Dumper.cdl
-- Created:	Fri Jun  3 09:43:20 1994
-- Author:	Christian CAILLET
--		<cky@sdsun2>
---Copyright:	 Matra Datavision 1994


class Dumper  from IGESSelect  inherits SessionDumper

    ---Purpose : Dumper from IGESSelect takes into account, for SessionFile, the
    --           classes defined in the package IGESSelect : Selections,
    --           Dispatches, Modifiers

uses Transient, AsciiString from TCollection, SessionFile

is

    Create returns mutable Dumper;
    ---Purpose : Creates a Dumper and puts it into the Library of Dumper

    WriteOwn (me; file : in out SessionFile; item : Transient) returns Boolean;
    ---Purpose : Write the Own Parameters of Types defined in package IGESSelect
    --           Returns True if <item> has been processed, False else

    ReadOwn  (me; file : in out SessionFile;
    	    type : AsciiString from TCollection; item : out mutable Transient)
    	returns Boolean;
    ---Purpose : Recognizes and Read Own Parameters for Types of package
    --           IGESSelect. Returns True if done and <item> created, False else

end Dumper;
