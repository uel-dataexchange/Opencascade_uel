-- File:	BRepAlgoAPI_Common.cdl
-- Created:	Thu Oct 14 18:25:52 1993
-- Author:	Remi LEQUETTE
--		<rle@phylox>
---Copyright:	 Matra Datavision 1993



class Common from BRepAlgoAPI inherits BooleanOperation from BRepAlgoAPI

	---Purpose: The class Common provides a
    	-- Boolean common operation on a pair of arguments (Boolean Intersection).
    	--  The class Common provides a framework for:
    	-- -           Defining the construction of a common shape;
    	-- -           Implementing the   building algorithm
    	-- -           Consulting the result.

uses
    Shape from TopoDS, 
    DSFiller from BOPTools

is
    Create (S1,S2 : Shape from TopoDS)  
    	returns Common from BRepAlgoAPI;  
	---Purpose: Constructs a common part for shapes aS1 and aS2 .
 
    Create (S1,S2 : Shape from TopoDS; 
    	    aDSF:DSFiller from BOPTools)  
    	returns Common from BRepAlgoAPI;
end Common;
--- Purpose: Constructs a common part for shapes aS1 and aS2 using aDSFiller
