-- File:        PlusMinusTolerance.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPlusMinusTolerance from RWStepShape

	---Purpose : Read & Write Module for PlusMinusTolerance

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PlusMinusTolerance from StepShape,
     EntityIterator from Interface

is

	Create returns RWPlusMinusTolerance;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PlusMinusTolerance from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : PlusMinusTolerance from StepShape);

	Share(me; ent : PlusMinusTolerance from StepShape; iter : in out EntityIterator);

end RWPlusMinusTolerance;
