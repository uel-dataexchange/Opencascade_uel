-- File:	BOPTools_Tools2D.cdl
-- Created:	Mon Apr  2 12:20:21 2001
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2001


class Tools2D from BOPTools 

	---Purpose: 
    	---  The class contains handy static functions 
	---  dealing with the topology 
uses 
    Vec  from gp, 
    Dir  from gp, 
    Vertex from TopoDS,
    Edge   from TopoDS, 
    Face   from TopoDS, 
     
    Curve from Geom2d,
    Curve from Geom, 
    ProjectedCurve from ProjLib

is   

    RemovePCurveForEdgeOnFace  (myclass; 
    	    	     aE:  Edge from TopoDS; 
                     aF:  Face from TopoDS); 
    	---Purpose: 
    	--- Remove P-Curve of the edge <aE> on the face <aF> 
    	---
    BuildPCurveForEdgeOnFace  (myclass; 
    	    	     aE:  Edge from TopoDS; 
                     aF:  Face from TopoDS); 
    	---Purpose: 
    	--- Compute P-Curve for the edge <aE> on the face <aF> 
    	---
    EdgeTangent     (myclass;  
			anE  : Edge from TopoDS; 
			aT   : Real from Standard; 
    	    	    	Tau  : out Vec  from gp) 
    	returns  Boolean from Standard; 
    	---Purpose: 
    	--- Compute tangent for the edge  <aE> [in 3D]  at parameter <aT> 
    	---
    FaceNormal      (myclass; 
                     aF:  Face from TopoDS; 
    	    	     U :  Real from Standard; 
                     V :  Real from Standard;  
    	    	     aN: out Vec  from gp); 
    	---Purpose: 
    	--- Compute normal for the face <aF> at parameters <U,V> 
    	--- of the corresp. surface. 
    	---
    PointOnSurface  (myclass; 
                     aE:  Edge from TopoDS; 
                     aF:  Face from TopoDS;  
    	    	     aT:  Real from Standard; 
                     U : out Real from Standard; 
                     V : out Real from Standard); 
    	---Purpose: 
    	--- Compute surface parameters <U,V> of the face <aF> 
    	--- for  the point from the edge <aE> at parameter <aT>.   
    	---
    CurveOnSurface  (myclass; 
                     aE:  Edge from TopoDS; 
                     aF:  Face from TopoDS; 
                     aC    : out Curve from Geom2d; 
                     aToler: out Real from Standard; 
    	    	     aTrim3d:Boolean from Standard); 
    	---Purpose:  
    	--- Get P-Curve <aC>  for the edge <aE> on surface <aF> . 
    	--- If the P-Curve does not exist, build  it using Make2D(). 
    	--- [aToler] - reached tolerance 
    	--- [aTrim3d] - trimming flag. 
    	---
    CurveOnSurface  (myclass; 
                     aE:  Edge from TopoDS; 
                     aF:  Face from TopoDS; 
                     aC    : out Curve from Geom2d; 
                     aFirst: out Real from Standard; 
                     aLast : out Real from Standard; 
                     aToler: out Real from Standard; 
    	    	     aTrim3d:Boolean from Standard); 
                      
    	---Purpose: 
    	--- Get P-Curve <aC>  for the edge <aE> on surface <aF> . 
    	--- If the P-Curve does not exist, build  it using Make2D(). 
    	--- [aFirst, aLast] - range of the P-Curve    
    	--- [aToler] - reached tolerance 
    	--- [aTrim3d] - trimming flag. 
    	---
    HasCurveOnSurface  (myclass;  
    	    	        aE:  Edge from TopoDS; 
                        aF:  Face from TopoDS; 
                        aC    : out Curve from Geom2d;
                        aFirst: out Real from Standard; 
                        aLast : out Real from Standard; 
                        aToler: out Real from Standard) 
    	returns  Boolean from Standard; 
    	---Purpose:  
    	--- Returns TRUE if the edge <aE>  has  P-Curve <aC>  	 
    	--- on surface <aF> .   
    	--- [aFirst, aLast] - range of the P-Curve    
    	--- [aToler] - reached tolerance 
    	--- If the P-Curve does not exist, aC.IsNull()=TRUE. 
    	---
    HasCurveOnSurface  (myclass;  
    	    	        aE:  Edge from TopoDS; 
                        aF:  Face from TopoDS) 
    	returns  Boolean from Standard;  
    	---Purpose:  
    	--- Returns TRUE if the edge <aE>  has  P-Curve <aC>  	 
    	--- on surface <aF> .   
    	--- If the P-Curve does not exist, aC.IsNull()=TRUE. 
    	---
    MakeCurveOnSurface	(myclass;  
    	    	        aE:  Edge from TopoDS; 
                        aF:  Face from TopoDS; 
                        aC    : out Curve from Geom2d;
                        aFirst: out Real from Standard; 
                        aLast : out Real from Standard; 
                        aToler: out Real from Standard; 
    	    	    	aTrim3d:Boolean from Standard);    	 
	 
    	---Purpose:   
    	--- Same  as   Make2D() 
    	---
    Make2D           (myclass;  
    	    	        aE:  Edge from TopoDS; 
                        aF:  Face from TopoDS; 
                        aC    : out Curve from Geom2d;
                        aFirst: out Real from Standard; 
                        aLast : out Real from Standard; 
                        aToler: out Real from Standard; 
    	    	    	aTrim3d:Boolean from Standard);    	
    	---Purpose:   
    	--- Make P-Curve <aC> for the edge <aE> on surface <aF> . 
    	--- [aFirst, aLast] - range of the P-Curve    
    	--- [aToler] - reached tolerance 
    	--- [aTrim3d] - trimming flag. 
    	---
    MakePCurveOnFace  (myclass;    
    	    	    	aF:  Face from TopoDS; 
    	    	    	C3D   :     Curve from Geom; 
			aC    : out Curve from Geom2d; 
			aToler: out Real from Standard) ;   
    	---Purpose:   
    	--- Make P-Curve <aC> for the 3D-curve <C3D> on surface <aF> . 
    	--- [aToler] - reached tolerance 
    	---
    MakePCurveOnFace  (myclass;    
    	    	    	aF:  Face from TopoDS; 
    	    	    	C3D   :     Curve from Geom;  
			aT1   :  Real from Standard;   
			aT2   :  Real from Standard;      
			aC    : out Curve from Geom2d; 
			aToler: out Real from Standard) ;  		
    	---Purpose:   
    	--- Make P-Curve <aC> for the 3D-curve <C3D> on surface <aF> .  
    	--- [aT1,  aT2] - range to build    
    	--- [aToler] - reached tolerance 
    	---
    AdjustPCurveOnFace  (myclass;    
    	    	    	aF    :  Face from TopoDS; 
    	    	    	C3D   :  Curve from Geom; 
			aC2D  :  Curve from Geom2d; 
			aC2DA : out Curve from Geom2d); 		 
    	---Purpose:   
    	--- Adjust P-Curve <aC2D> (3D-curve <C3D>) on surface <aF> .  
    	---
    AdjustPCurveOnFace  (myclass;    
    	    	    	aF    :  Face from TopoDS; 
			aT1   :  Real from Standard;   
			aT2   :  Real from Standard;   
			aC2D  :  Curve from Geom2d; 
			aC2DA : out Curve from Geom2d); 
    	---Purpose:   
    	--- Adjust P-Curve <aC2D> (3D-curve <C3D>) on surface <aF> .  
    	--- [aT1,  aT2] - range to adjust 
    	---
    MakePCurveOfType  (myclass;    
    		       PC  : ProjectedCurve from ProjLib; 
    	    	       aC  : out Curve from Geom2d);	 
    	---Purpose:   
    	--- Make empty  P-Curve <aC> of relevant to <PC> type  
    	---
    TangentOnEdge    (myclass;  
    	    	    	aParm: Real from Standard; 
			anE  : Edge from TopoDS;  
			aTang: out Vec  from gp) 
    	returns  Boolean from Standard; 
    	---Purpose:   
    	--- Compute tangent for the edge <anE> at parameter <aParm>        
    	---
    TangentOnEdge    (myclass;  
			anE  : Edge from TopoDS;  
			aDTang: out Dir  from gp) 
    	returns  Boolean from Standard;  
    	---Purpose:   
    	--- Compute tangent for the edge <anE> at arbitrary intermediate parameter.        
    	---
    TangentOnVertex  (myclass;  
    	    	    	aVF  : Vertex from TopoDS; 
    	    	    	aVL  : Vertex from TopoDS; 
			anE  : Edge from TopoDS;  
			aTang: out  Vec  from gp) 
    	returns  Boolean from Standard;  
    	---Purpose:   
    	--- Compute tangent for the vertex point <aVF> for the edge <anE>. 
    	--- <aVL> is opposite vertex of the edge        
    	---
    EdgeBounds        (myclass; 
    	    	    	 anE  : Edge from TopoDS;   
			 aFirst: out Real from Standard; 
                         aLast : out Real from Standard); 
    	---Purpose:   
    	--- Returns parametric range for the edge <anE>. 
    	---
    IntermediatePoint (myclass; 
    	    	    	 aFirst: Real from Standard; 
                         aLast : Real from Standard) 
    	returns  Real from Standard; 
    	---Purpose:   
    	--- Compute intermediate  value in  between [aFirst, aLast] . 
    	---
    IntermediatePoint	(myclass;  
    	    	    	  anE  : Edge from TopoDS) 
	returns  Real from Standard;
    	---Purpose:   
    	--- Compute intermediate value of parameter for the edge <anE>. 
    	---

end Tools2D;
