-- File:	StepBasic_PhysicallyModeledProductDefinition.cdl
-- Created:	Tue Jun 30 15:58:33 1998
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1998


class PhysicallyModeledProductDefinition  from StepBasic
    inherits ProductDefinition  from StepBasic

uses
     HAsciiString from TCollection

is

    Create returns PhysicallyModeledProductDefinition;

end PhysicallyModeledProductDefinition;
