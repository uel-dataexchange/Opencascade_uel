-- File:	IGESDimen_ToolCenterLine.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolCenterLine  from IGESDimen

    ---Purpose : Tool to work on a CenterLine. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses CenterLine from IGESDimen,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolCenterLine;
    ---Purpose : Returns a ToolCenterLine, ready to work


    ReadOwnParams (me; ent : mutable CenterLine;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : CenterLine;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : CenterLine;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a CenterLine <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable CenterLine) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a CenterLine
    --           (LineFont forced to Rank = 1, DataType forced to 1)

    DirChecker (me; ent : CenterLine) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : CenterLine;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : CenterLine; entto : mutable CenterLine;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : CenterLine;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolCenterLine;
