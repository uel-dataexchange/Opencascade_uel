-- File:	Transfer_ActorOfFinderProcess.cdl
-- Created:	Wed Sep  4 17:44:43 1996
-- Author:	Christian CAILLET
--		<cky@fidox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996


class ActorOfFinderProcess  from Transfer  inherits ActorOfProcessForFinder

    ---Purpose : The original class was renamed. Compatibility only
    --         
    --         ModeTrans : a simple way of transmitting a transfer mode from
    --         a user. To be interpreted for each norm

uses Finder, FinderProcess, ProcessForFinder, Binder

is

    Create  returns mutable ActorOfFinderProcess;

    ModeTrans (me : mutable) returns Integer;
    ---Purpose : Returns the Transfer Mode, modifiable
    ---C++ : return &

    Transferring (me : mutable; start : Finder; TP : mutable ProcessForFinder)
        returns mutable Binder  is redefined;
    -- calls the one below

    Transfer (me : mutable; start : Finder; TP : mutable FinderProcess)
        returns mutable Binder  is virtual;
    -- default calls TransferTransient if <start> is a TransientMapper,
    -- i.e. does nothing, to be redefined

    TransferTransient (me : mutable; start : Transient;
    	    	       TP : mutable FinderProcess)
	returns mutable Transient  is virtual;
    -- default does nothing, can be redefined
    -- usefull when a result is Transient, simpler to define than Transfer with
    -- a Finder

fields

    themodetrans : Integer  is protected;

end ActorOfFinderProcess;
