-- File:	IGESSelect_ComputeStatus.cdl
-- Created:	Wed Jun  1 16:18:06 1994
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1994


class ComputeStatus  from IGESSelect  inherits ModelModifier from IGESSelect

    ---Purpose : Computes Status of IGES Entities for a whole IGESModel.
    --           This concerns SubordinateStatus and UseFlag, which must have
    --           some definite values according the way they are referenced.
    --           (see definitions of Logical use, Physical use, etc...)
    --           
    --           Works by calling a BasicEditor from IGESData. Works on the
    --           whole produced (target) model, because computation is global.

uses AsciiString from TCollection,
     IGESModel, CopyTool, ContextModif

is

    Create returns mutable ComputeStatus;
    ---Purpose : Creates an ComputeStatus, which uses the system Date


    Performing (me; ctx : in out ContextModif;
    	        target  : mutable IGESModel;
                TC      : in out CopyTool);
    ---Purpose : Specific action : it first evaluates the required values for
    --           Subordinate Status and Use Flag (in Directory Part of each
    --           IGES Entity). Then it corrects them, for the whole target.
    --           Works with a Protocol. Implementation uses BasicEditor

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text which is
    --           "Compute Subordinate Status and Use Flag"

end ComputeStatus;
