-- File:	PDataStd_ExtStringArray_1.cdl
-- Created:	Thu Mar 27 17:09:57 2008
-- Author:	Sergey ZARITCHNY
--		<sergey.zaritchny@opencascade.com>
---Copyright:	Open CasCade SA 2008 

class ExtStringArray_1 from PDataStd inherits Attribute from PDF

	---Purpose: Persistence

uses  HExtendedString          from PCollection,
      HArray1OfExtendedString  from PColStd
     
     
is

    Create returns mutable ExtStringArray_1 from PDataStd;

    Init(me : mutable; lower, upper : Integer from Standard);

    SetValue(me: mutable; Index : Integer from Standard; Value : HExtendedString from PCollection);
    
    Value(me;  Index : Integer from Standard) returns HExtendedString from PCollection;
   
    Lower (me) returns Integer from Standard;      

    Upper (me) returns Integer from Standard;   
     
    SetDelta(me : mutable; delta : Boolean from Standard); 
     
    GetDelta(me) returns Boolean from Standard;
     
fields
    myValue     :  HArray1OfExtendedString from PColStd;
    myDelta  : Boolean from Standard;

end ExtStringArray_1;



