-- File:	StepData_Plex.cdl
-- Created:	Fri May  9 16:35:59 1997
-- Author:	Christian CAILLET
--		<cky@heliox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


class Plex  from StepData    inherits Described  from StepData

    ---Purpose : A Plex (for Complex) Entity is defined as a list of Simple
    --           Members ("external mapping")
    --           The types of these members must be in alphabetic order

uses CString,
     SequenceOfTransient from TColStd,
     HSequenceOfAsciiString from TColStd,
     Check from Interface,  EntityIterator from Interface,
     ECDescr from StepData, Simple from StepData, Field from StepData

raises InterfaceMismatch

is

    Create (descr : ECDescr) returns mutable Plex;
    ---Purpose : Creates a Plex (empty). The complete creation is made by the
    --           ECDescr itself, by calling Add

    Add (me : mutable; member : Simple);
    ---Purpose : Adds a member to <me>

    ECDescr (me) returns ECDescr;
    ---Purpose : Returns the Description as for a Plex

    	--  inherited

    IsComplex (me) returns Boolean;
    ---Purpose : Returns False


    Matches (me; steptype : CString) returns Boolean;
    ---Purpose : Tells if a step type is matched by <me>
    --           For a Simple Entity : own type or super type
    --           For a Complex Entity : one of the members

    As (me; steptype : CString) returns mutable Simple;
    ---Purpose : Returns a Simple Entity which matches with a Type in <me> :
    --           For a Simple Entity : me if it matches, else a null handle
    --           For a Complex Entity : the member which matches, else null

    HasField (me; name : CString) returns Boolean;
    ---Purpose : Tells if a Field brings a given name

    Field (me; name : CString) returns Field
    ---Purpose : Returns a Field from its name; read-only
    	raises InterfaceMismatch;
    --           raises if no Field for <name>
    ---C++ : return const &

    CField (me : mutable; name : CString) returns Field
    ---Purpose : Returns a Field from its name; read or write
    	raises InterfaceMismatch;
    --           raises if no Field for <name>
    ---C++ : return &

    	-- more specific

    NbMembers (me) returns Integer;
    ---Purpose : Returns the count of simple members

    Member (me; num : Integer) returns Simple;
    ---Purpose : Returns a simple member from its rank

    TypeList (me) returns HSequenceOfAsciiString;
    ---Purpose : Returns the actual list of members types

    	--

    Check  (me; ach  : in out Check from Interface);
    ---Purpose : Fills a Check by using its Description

    Shared (me; list : in out EntityIterator from Interface);
    ---Purpose : Fills an EntityIterator with entities shared by <me>

fields

    themembers : SequenceOfTransient;

end Plex;
