-- File:	IGESBasic_SpecificModule.cdl
-- Created:	Tue Sep  7 11:14:37 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class SpecificModule  from IGESBasic  inherits  SpecificModule from IGESData

    ---Purpose : Defines Services attached to IGES Entities :
    --           Dump & OwnCorrect, for IGESBasic

uses IGESEntity, IGESDumper,
     Messenger from Message

is

    Create returns mutable SpecificModule from IGESBasic;
    ---Purpose : Creates a SpecificModule from IGESBasic & puts it into SpecificLib

    OwnDump (me; CN : Integer; ent : IGESEntity;
    	      dumper : IGESDumper;  S : Messenger from Message; own : Integer);
    ---Purpose : Specific Dump (own parameters) for IGESBasic

    OwnCorrect (me; CN : Integer; ent : mutable IGESEntity)
    	returns Boolean  is redefined;
    ---Purpose : Performs non-ambiguous Corrections on Entities which support
    --           them (AssocGroupType,Hierarchy,Name,SingleParent)

end SpecificModule;
