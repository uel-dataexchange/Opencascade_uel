-- File:	IGESAppli_ToolRegionRestriction.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolRegionRestriction  from IGESAppli

    ---Purpose : Tool to work on a RegionRestriction. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses RegionRestriction from IGESAppli,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolRegionRestriction;
    ---Purpose : Returns a ToolRegionRestriction, ready to work


    ReadOwnParams (me; ent : mutable RegionRestriction;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : RegionRestriction;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : RegionRestriction;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a RegionRestriction <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable RegionRestriction) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a RegionRestriction
    --           (NbPropertyValues forced to 3, Level cleared if Subordinate != 0)

    DirChecker (me; ent : RegionRestriction) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : RegionRestriction;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : RegionRestriction; entto : mutable RegionRestriction;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : RegionRestriction;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolRegionRestriction;
