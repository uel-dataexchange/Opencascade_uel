-- File:	IGESGeom_ToolBSplineSurface.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolBSplineSurface  from IGESGeom

    ---Purpose : Tool to work on a BSplineSurface. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses BSplineSurface from IGESGeom,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolBSplineSurface;
    ---Purpose : Returns a ToolBSplineSurface, ready to work


    ReadOwnParams (me; ent : mutable BSplineSurface;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : BSplineSurface;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : BSplineSurface;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a BSplineSurface <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : BSplineSurface) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : BSplineSurface;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : BSplineSurface; entto : mutable BSplineSurface;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : BSplineSurface;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolBSplineSurface;
