-- File:	BinMDataStd_ExtStringArrayDriver.cdl
-- Created:	Tue Aug 24 17:19:27 2004
-- Author:	Pavel TELKOV
--		<ptv@valenox>
---Copyright:	 Matra Datavision 2004

class ExtStringArrayDriver from BinMDataStd inherits ADriver from BinMDF

        ---Purpose: Array of extended string attribute Driver.

uses
    MessageDriver    from CDM,
    SRelocationTable from BinObjMgt,
    RRelocationTable from BinObjMgt,
    Persistent       from BinObjMgt,
    Attribute        from TDF

is
    Create (theMessageDriver:MessageDriver from CDM)
        returns mutable ExtStringArrayDriver from BinMDataStd;

    NewEmpty (me)  returns mutable Attribute from TDF
    	is redefined;

    Paste(me; Source     : Persistent from BinObjMgt;
              Target     : mutable Attribute from TDF;
              RelocTable : out RRelocationTable from BinObjMgt)
        returns Boolean from Standard is redefined;

    Paste(me; Source     : Attribute from TDF;
              Target     : in out Persistent from BinObjMgt;
              RelocTable : out SRelocationTable from BinObjMgt)
    	is redefined;

end ExtStringArrayDriver;
