-- File:        SurfaceReplica.cdl
-- Created:     Mon Dec  4 12:02:31 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWSurfaceReplica from RWStepGeom

	---Purpose : Read & Write Module for SurfaceReplica

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     SurfaceReplica from StepGeom,
     EntityIterator from Interface

is

	Create returns RWSurfaceReplica;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable SurfaceReplica from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : SurfaceReplica from StepGeom);

	Share(me; ent : SurfaceReplica from StepGeom; iter : in out EntityIterator);

end RWSurfaceReplica;
