-- File:        PresentationLayerUsage.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPresentationLayerUsage from RWStepVisual

	---Purpose : Read & Write Module for PresentationLayerUsage

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PresentationLayerUsage from StepVisual,
     EntityIterator from Interface

is

	Create returns RWPresentationLayerUsage;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PresentationLayerUsage from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : PresentationLayerUsage from StepVisual);

	Share(me; ent : PresentationLayerUsage from StepVisual; iter : in out EntityIterator);

end RWPresentationLayerUsage;
