-- File:	StepToGeom_MakeTrimmedCurve.cdl
-- Created:	Fri Nov  4 10:28:03 1994
-- Author:	Frederic MAUPAS
---Copyright:	 Matra Datavision 1994

class MakeTrimmedCurve2d from StepToGeom

    ---Purpose: This class implements the mapping between classes 
    --          class TrimmedCurve from StepGeom which
    --          describes a Trimmed Curve from prostep and TrimmedCurve from 
    --          Geom. 
  
uses BSplineCurve from Geom2d,
     TrimmedCurve from StepGeom

is 

    Convert ( myclass; SC : TrimmedCurve from StepGeom;
                       CC : out BSplineCurve from Geom2d )
    returns Boolean from Standard;

end MakeTrimmedCurve2d;
