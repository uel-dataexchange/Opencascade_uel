-- File:	IGESAppli_ToolFiniteElement.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolFiniteElement  from IGESAppli

    ---Purpose : Tool to work on a FiniteElement. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses FiniteElement from IGESAppli,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolFiniteElement;
    ---Purpose : Returns a ToolFiniteElement, ready to work


    ReadOwnParams (me; ent : mutable FiniteElement;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : FiniteElement;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : FiniteElement;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a FiniteElement <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : FiniteElement) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : FiniteElement;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : FiniteElement; entto : mutable FiniteElement;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : FiniteElement;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolFiniteElement;
