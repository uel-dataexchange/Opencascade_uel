-- File:	StepData_FileProtocol.cdl
-- Created:	Fri Jul 23 10:13:04 1993
-- Author:	Christian CAILLET
--		<cky@meteox>
---Copyright:	 Matra Datavision 1993


class FileProtocol  from StepData  inherits Protocol from StepData

    ---Purpose : A FileProtocol is defined as the addition of several already
    --           existing Protocols. It corresponds to the definition of a
    --           SchemaName with several Names, each one being attached to a
    --           specific Protocol. Thus, a File defined with a compound Schema
    --           is processed as any other one, once built the equivalent
    --           compound Protocol, a FileProtocol

uses Type, CString, SequenceOfTransient,
     Graph from Interface, Check from Interface,
     Protocol from Interface, Protocol from StepData

is

    Create returns mutable FileProtocol;
    ---Purpose : Creates an empty FileProtocol

    Add (me : mutable; protocol : Protocol from StepData);
    ---Purpose : Adds a Protocol to the definition list of the FileProtocol
    --           But ensures that each class of Protocol is present only once
    --           in this list

    NbResources (me) returns Integer  is redefined;
    ---Purpose : Gives the count of Protocols used as Resource (can be zero)
    --           i.e. the count of Protocol recorded by calling the method Add

    Resource (me; num : Integer) returns Protocol from Interface  is redefined;
    ---Purpose : Returns a Resource, given a rank. Here, rank of calling Add

    TypeNumber (me; atype : any Type) returns Integer  is redefined;
    ---Purpose : Returns a Case Number, specific of each recognized Type
    --           Here, NO Type at all is recognized properly : all Types are
    --           recognized by the resources

    GlobalCheck (me; G : Graph; ach : in out Check)
    	returns Boolean  is redefined;
    ---Purpose : Calls GlobalCheck for each of its recorded ressources

    	-- --    Specific for StepData    -- --

    SchemaName (me) returns CString  is redefined;
    ---Purpose : Returns the Schema Name attached to each class of Protocol
    --           To be redefined by each sub-class
    --           Here, SchemaName returns "" (empty String)
    -- was C++ : return const

fields

    thecomps : SequenceOfTransient;

end FileProtocol;
