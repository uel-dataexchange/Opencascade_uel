-- File:	IGESDefs_SpecificModule.cdl
-- Created:	Tue Sep  7 11:14:37 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class SpecificModule  from IGESDefs  inherits  SpecificModule from IGESData

    ---Purpose : Defines Services attached to IGES Entities : Dump, for IGESDefs

uses Messenger from Message, IGESEntity, IGESDumper

is

    Create returns mutable SpecificModule from IGESDefs;
    ---Purpose : Creates a SpecificModule from IGESDefs & puts it into SpecificLib

    OwnDump (me; CN : Integer; ent : IGESEntity;
    	      dumper : IGESDumper;  S : Messenger from Message; own : Integer);
    ---Purpose : Specific Dump (own parameters) for IGESDefs

end SpecificModule;
