-- File:	StepElement_Curve3dElementDescriptor.cdl
-- Created:	Thu Dec 12 17:28:59 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class Curve3dElementDescriptor from StepElement
inherits ElementDescriptor from StepElement

    ---Purpose: Representation of STEP entity Curve3dElementDescriptor

uses
    ElementOrder from StepElement,
    HAsciiString from TCollection,
    HArray1OfHSequenceOfCurveElementPurposeMember from StepElement

is
    Create returns Curve3dElementDescriptor from StepElement;
	---Purpose: Empty constructor

    Init (me: mutable; aElementDescriptor_TopologyOrder: ElementOrder from StepElement;
                       aElementDescriptor_Description: HAsciiString from TCollection;
                       aPurpose: HArray1OfHSequenceOfCurveElementPurposeMember from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    Purpose (me) returns HArray1OfHSequenceOfCurveElementPurposeMember from StepElement;
	---Purpose: Returns field Purpose
    SetPurpose (me: mutable; Purpose: HArray1OfHSequenceOfCurveElementPurposeMember from StepElement);
	---Purpose: Set field Purpose

fields
    
    thePurpose: HArray1OfHSequenceOfCurveElementPurposeMember from StepElement;

end Curve3dElementDescriptor;
