-- File:	RWStepShape_RWSeamEdge.cdl
-- Created:	Fri Jan  4 17:42:44 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWSeamEdge from RWStepShape

    ---Purpose: Read & Write tool for SeamEdge

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    SeamEdge from StepShape

is
    Create returns RWSeamEdge from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : SeamEdge from StepShape);
	---Purpose: Reads SeamEdge

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: SeamEdge from StepShape);
	---Purpose: Writes SeamEdge

    Share (me; ent : SeamEdge from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWSeamEdge;
