-- File:        CameraModelD3.cdl
-- Created:     Fri Dec  1 11:11:15 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class CameraModelD3 from StepVisual 

inherits CameraModel from StepVisual 

uses

	Axis2Placement3d from StepGeom, 
	ViewVolume from StepVisual, 
	HAsciiString from TCollection
is

	Create returns mutable CameraModelD3;
	---Purpose: Returns a CameraModelD3


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aViewReferenceSystem : mutable Axis2Placement3d from StepGeom;
	      aPerspectiveOfVolume : mutable ViewVolume from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetViewReferenceSystem(me : mutable; aViewReferenceSystem : mutable Axis2Placement3d);
	ViewReferenceSystem (me) returns mutable Axis2Placement3d;
	SetPerspectiveOfVolume(me : mutable; aPerspectiveOfVolume : mutable ViewVolume);
	PerspectiveOfVolume (me) returns mutable ViewVolume;

fields

	viewReferenceSystem : Axis2Placement3d from StepGeom;
	perspectiveOfVolume : ViewVolume from StepVisual;

end CameraModelD3;
