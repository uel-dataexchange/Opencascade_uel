-- File:	IGESSolid_ToolSolidAssembly.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolSolidAssembly  from IGESSolid

    ---Purpose : Tool to work on a SolidAssembly. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses SolidAssembly from IGESSolid,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolSolidAssembly;
    ---Purpose : Returns a ToolSolidAssembly, ready to work


    ReadOwnParams (me; ent : mutable SolidAssembly;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : SolidAssembly;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : SolidAssembly;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a SolidAssembly <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : SolidAssembly) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : SolidAssembly;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : SolidAssembly; entto : mutable SolidAssembly;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : SolidAssembly;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolSolidAssembly;
