-- File:	TCompSolid1.cdl
-- Created:	Mon Dec 17 11:18:44 1990
-- Author:	Remi Lequette
--		<rle@topsn3>
---Copyright:	 Matra Datavision 1990, 1992



class TCompSolid1 from PTopoDS inherits TShape1 from PTopoDS

	---Purpose: A  topological Composite  Solid1 shape.

uses
    ShapeEnum from TopAbs

is
    Create returns mutable TCompSolid1 from PTopoDS;
	---Purpose: The new  TCompSolid11 is empty.
    ---Level: Internal 
    	
    ShapeType(me) returns ShapeEnum from TopAbs;
    ---Level: Internal 

end TCompSolid1;
