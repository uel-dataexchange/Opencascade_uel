-- File:	BRepBuilderAPI_Transform.cdl
-- Created:	Fri Dec  9 09:02:17 1994
-- Author:	Jacques GOUSSARD
--		<jag@topsn2>
---Copyright:	 Matra Datavision 1994


class Transform from BRepBuilderAPI inherits ModifyShape from BRepBuilderAPI

	---Purpose: Geometric transformation on a shape.
    	-- The transformation to be applied is defined as a
    	-- gp_Trsf transformation, i.e. a transformation which does
    	-- not modify the underlying geometry of shapes.
    	-- The transformation is applied to:
    	-- -   all curves which support edges of a shape, and
    	-- -   all surfaces which support its faces.
    	-- A Transform object provides a framework for:
    	-- -   defining the geometric transformation to be applied,
    	-- -   implementing the transformation algorithm, and
    	-- -   consulting the results.
    
uses 
    Trsf              from gp,
    Location          from TopLoc,
    Shape             from TopoDS,
    Face              from TopoDS,
    ShapeModification from BRepBuilderAPI,
    ListOfShape       from TopTools

raises
 NoSuchObject from Standard    
is

    Create(T: Trsf from gp)
        
    	returns Transform from BRepBuilderAPI;
	---Purpose:  Constructs a framework for applying the geometric
    	-- transformation T to a shape. Use the function Perform
    	-- to define the shape to transform.


    Create(S: Shape from TopoDS; T: Trsf from gp; 
           Copy: Boolean from Standard  =  Standard_False)

    	returns Transform from BRepBuilderAPI;
	---Purpose: Creates a transformation from the gp_Trsf <T>, and
	--          applies it to the shape <S>. If the transformation
	--          is  direct   and isometric (determinant  =  1) and
	--          <Copy> =  Standard_False,  the resulting shape  is
	--          <S> on   which  a  new  location has    been  set.
	--          Otherwise,  the   transformation is applied   on a
	--          duplication of <S>.


    Perform(me: in out; S   : Shape   from TopoDS; 
                        Copy: Boolean from Standard  =  Standard_False)

	---Purpose: pplies the geometric transformation defined at the
    	-- time of construction of this framework to the shape S.
    	-- - If the transformation T is direct and isometric, in
    	-- other words, if the determinant of the vectorial part
    	-- of T is equal to 1., and if Copy equals false (the
    	-- default value), the resulting shape is the same as
    	-- the original but with a new location assigned to it.
    	-- -   In all other cases, the transformation is applied to a duplicate of S.
    	-- Use the function Shape to access the result.
    	-- Note: this framework can be reused to apply the same
    	-- geometric transformation to other shapes. You only
    	-- need to specify them by calling the function Perform again.

    	is static;

    ModifiedShape(me; S: Shape from TopoDS)
    	returns Shape from TopoDS
	---Purpose: Returns the modified shape corresponding to <S>.
	---C++: return const&
	raises NoSuchObject from Standard
               -- if S is not the initial shape or a sub-shape
               -- of the initial shape.
    is redefined virtual;

    Modified (me: in out; S : Shape from TopoDS)
    	---Purpose: Returns the list  of shapes modified from the shape
    	--          <S>. 
        ---C++: return const & 
        ---Level: Public
    returns ListOfShape from TopTools
    is redefined virtual;


fields

    myTrsf     : Trsf     from gp;
    myLocation : Location from TopLoc;
    myUseModif : Boolean  from Standard;
    
end Transform;
