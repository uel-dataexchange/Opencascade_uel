-- File:	StepShape_ConnectedEdgeSet.cdl
-- Created:	Fri Dec 28 16:02:00 2001 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class ConnectedEdgeSet from StepShape
inherits TopologicalRepresentationItem from StepShape

    ---Purpose: Representation of STEP entity ConnectedEdgeSet

uses
    HAsciiString from TCollection,
    HArray1OfEdge from StepShape

is
    Create returns ConnectedEdgeSet from StepShape;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aCesEdges: HArray1OfEdge from StepShape);
	---Purpose: Initialize all fields (own and inherited)

    CesEdges (me) returns HArray1OfEdge from StepShape;
	---Purpose: Returns field CesEdges
    SetCesEdges (me: mutable; CesEdges: HArray1OfEdge from StepShape);
	---Purpose: Set field CesEdges

fields
    theCesEdges: HArray1OfEdge from StepShape;

end ConnectedEdgeSet;
