-- File:	StepShape_ShapeRepresentationWithParameters.cdl
-- Created:	Wed Jun  4 13:34:33 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class ShapeRepresentationWithParameters from StepShape
inherits ShapeRepresentation from StepShape

    ---Purpose: Representation of STEP entity ShapeRepresentationWithParameters

uses
    HAsciiString from TCollection,
    HArray1OfRepresentationItem from StepRepr,
    RepresentationContext from StepRepr

is
    Create returns ShapeRepresentationWithParameters from StepShape;
	---Purpose: Empty constructor

end ShapeRepresentationWithParameters;
