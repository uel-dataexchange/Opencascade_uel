-- File:	MNaming_NamedShapeRetrievalDriver.cdl
-- Created:	Fri Apr 11 16:03:36 1997
-- Author:	VAUTHIER Jean-Claude
---Copyright:	 Matra Datavision 1997


class NamedShapeRetrievalDriver from MNaming inherits ARDriver from MDF

	---Purpose: 

uses
    RRelocationTable from MDF,
    Attribute        from PDF,
    Attribute        from TDF, 
    MessageDriver    from CDM


is


    Create(theMessageDriver : MessageDriver from CDM) -- Version 0
    returns mutable NamedShapeRetrievalDriver from MNaming;

    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type NamedShape from PNaming.

    NewEmpty (me)
    returns mutable Attribute from TDF;


    Paste(me;
    	  Source     :          Attribute        from PDF;
    	  Target     : mutable  Attribute        from TDF;
    	  RelocTable :          RRelocationTable from MDF);


end NamedShapeRetrievalDriver;
