-- File:	RWStepElement_RWAnalysisItemWithinRepresentation.cdl
-- Created:	Thu Dec 12 17:28:59 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWAnalysisItemWithinRepresentation from RWStepElement

    ---Purpose: Read & Write tool for AnalysisItemWithinRepresentation

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    AnalysisItemWithinRepresentation from StepElement

is
    Create returns RWAnalysisItemWithinRepresentation from RWStepElement;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : AnalysisItemWithinRepresentation from StepElement);
	---Purpose: Reads AnalysisItemWithinRepresentation

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: AnalysisItemWithinRepresentation from StepElement);
	---Purpose: Writes AnalysisItemWithinRepresentation

    Share (me; ent : AnalysisItemWithinRepresentation from StepElement;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWAnalysisItemWithinRepresentation;
