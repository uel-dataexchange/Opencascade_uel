-- File:	RWStepDimTol.cdl
-- Created:	Wed Jun  4 12:04:38 2003
-- Author:	Galina KULIKOVA
--		<gka@zamox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 2003


package RWStepDimTol 

	---Purpose: Packsge contains tools for parsing and formatting GD&T entities.

    uses
    	TCollection,
    	RWStepRepr, 
    	RWStepShape,
    	RWStepVisual,
    	RWStepBasic,
    	TColStd,
	StepData,
    	Interface, 
	StepDimTol,
    	MMgt

    is
    	class RWAngularityTolerance;
    	class RWCircularRunoutTolerance;
    	class RWConcentricityTolerance;
    	class RWCylindricityTolerance;
    	class RWCoaxialityTolerance;
    	class RWFlatnessTolerance;
    	class RWLineProfileTolerance;
    	class RWParallelismTolerance;
    	class RWPerpendicularityTolerance;
    	class RWPositionTolerance;
    	class RWRoundnessTolerance;
    	class RWStraightnessTolerance;
    	class RWSurfaceProfileTolerance;
    	class RWSymmetryTolerance;
    	class RWTotalRunoutTolerance;
    
    	class RWGeometricTolerance;
    	class RWGeometricToleranceRelationship;
    	class RWGeometricToleranceWithDatumReference;
    	class RWModifiedGeometricTolerance;
     
    	class RWDatum;
    	class RWDatumFeature;
    	class RWDatumReference;
    	class RWCommonDatum;
    	class RWDatumTarget;
    	class RWPlacedDatumTargetFeature;
    	
	class RWGeoTolAndGeoTolWthDatRefAndModGeoTolAndPosTol;


end RWStepDimTol;
