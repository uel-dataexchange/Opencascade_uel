-- File:	StepShape_Subedge.cdl
-- Created:	Fri Jan  4 17:42:45 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class Subedge from StepShape
inherits Edge from StepShape

    ---Purpose: Representation of STEP entity Subedge

uses
    HAsciiString from TCollection,
    Vertex from StepShape,
    Edge from StepShape

is
    Create returns Subedge from StepShape;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentationItem_Name: HAsciiString from TCollection;
                       aEdge_EdgeStart: Vertex from StepShape;
                       aEdge_EdgeEnd: Vertex from StepShape;
                       aParentEdge: Edge from StepShape);
	---Purpose: Initialize all fields (own and inherited)

    ParentEdge (me) returns Edge from StepShape;
	---Purpose: Returns field ParentEdge
    SetParentEdge (me: mutable; ParentEdge: Edge from StepShape);
	---Purpose: Set field ParentEdge

fields
    theParentEdge: Edge from StepShape;

end Subedge;
