
-- File:        Graphic2d_Drawer.cdl
-- Created:     Thu Jul  8 09:27:11 1993
-- Author:      Jean Louis FRENKEL
--              <jlf@stylox>
---
-- Modified : DCB 22-07-98
-- Reason   : Using pointers to drivers instead of handles
--
--            SAV 14/11/01 added MapMarkersFromTo(). operates with arrays.
--            
---Copyright:    Matra Datavision 1993

class Drawer from Graphic2d inherits Transient from Standard

        ---Version:

        ---Purpose: A Drawer groups all conversion methods.
        ---Level: Internal

        ---Keywords:
        ---Warning:
        ---References:

uses
        ShortReal               from Standard,
        File                    from OSD,
        Factor                  from Quantity,
        Driver                  from Aspect,
        DriverPtr               from Aspect,
        WindowDriver            from Aspect,
        WindowDriverPtr         from Aspect,
        PlotterDriver           from PlotMgt,
        PlotterDriverPtr        from PlotMgt,
        TypeOfDeflection        from Aspect,
        TypeOfText              from Aspect,
        Array1OfShortReal       from TShort,
        ExtendedString          from TCollection,
	HArray1OfShortReal      from TShort

raises
        DrawerDefinitionError   from Graphic2d

is
        -------------------------
        -- Category: Constructors
        -------------------------

        Create
        returns mutable Drawer from Graphic2d;
        ---Level: Internal
        ---Purpose: A drawer is :
        --      - a driver
        --      - a "map from" and a "map to"
        --      - attributes
        ---Category: Constructors

        -----------------------------------------
        -- Category: Methods to modify the driver
        -----------------------------------------

        SetDriver (me: mutable; aDriver: Driver from Aspect)
                is static;
        ---Level: Internal
        ---Purpose: Associates the driver <ADriver> to the drawer <me>.
        ---Category: Methods to modify the driver

        Driver (me)
                returns Driver from Aspect
        ---Level: Internal
        ---Purpose: Returns the associated driver.
        --  Warning: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;

        IsWindowDriver (me) 
                returns Boolean from Standard;
        ---Level: Internal
        ---Purpose: Returns TRUE if the driver is a window driver.
        ---Category: Inquiry method.

        WindowDriver (me)
                returns WindowDriver from Aspect
        ---Level: Internal
        ---Purpose: Returns the associated window driver.
        --  Warning: Raises DrawerDefinitionError if the
        --          associated driver is not defined or is not a WindowDriver.
        raises DrawerDefinitionError from Graphic2d is static;

        IsPlotterDriver (me) 
                returns Boolean from Standard;
        ---Level: Internal
        ---Purpose: Returns TRUE if the driver is a plotter driver.
        ---Category: Inquiry method.

        PlotterDriver (me)
                returns PlotterDriver from PlotMgt
        ---Level: Internal
        ---Purpose: Returns the associated plotter driver.
        --  Warning: Raises DrawerDefinitionError if the
        --          associated driver is not defined or is not a PlotterDriver
        raises DrawerDefinitionError from Graphic2d is static;

        ----------------------------------------------------
        -- Category: Methods to modify the chordal deviation
        ----------------------------------------------------

        ----------------------------------------------------------
        -- Summary of chordal deviation                         --
        --                                                      --
        -- Specify a chordal deviation that is smaller than the --
        -- workstation pixel size will not improve the display, --
        -- but will slow the drawing.                           --
        --                                                      --
        ----------------------------------------------------------

        SetDrawPrecision (me: mutable; aPrecision: Real from Standard;
                aCoefficient: Real from Standard;
                aType: TypeOfDeflection from Aspect)
                is static;
        ---Level: Internal
        ---Purpose: Sets the chordal deviation.
        --          <aPrecision> is the chordal deviation when the type of
        --          deflection is Aspect_TOD_ABSOLUTE.
        --          <aCoefficient> is used when when the type of
        --          deflection is Aspect_TOD_RELATIVE.
        --      TypeOfDeflection is :
        --              Aspect_TOD_RELATIVE
        --              Aspect_TOD_ABSOLUTE
        --      TypeOfDeflection defines if the maximal chordal deviation
        --      used when drawing an object is absolute or relative to the
        --      size of the object.
        --  Warning: Specify a chordal deviation that is smaller than the
        --          workstation pixel size will not improve the display,
        --          but will slow the drawing.

        DrawPrecision (me; aPrecision: out ShortReal from Standard;
                aCoefficient: out ShortReal from Standard;
                aType: out TypeOfDeflection from Aspect)
                is static;
        ---Level: Internal
        ---Purpose: Returns the chordal deviation.

        SetTextPrecision (me: mutable; aPrecision: ShortReal from Standard)
                is static;
        ---Level: Internal
        ---Purpose: Sets the Text precision in METER
        -- Any text is displayed only if his height is greater than
        --the text precision or replaced by a bounding box in the other case.

        TextPrecision (me) returns ShortReal from Standard
                is static;
        ---Level: Internal
        ---Purpose: Returns the Text precision in METER.

        ---------------------------------------------
        -- Category: Methods to modify the 2D viewing
        ---------------------------------------------

        SetValues (me: mutable; XF, YF, SF, XT, YT, ST, ZF: Real from Standard)
                is static;
        ---Level: Internal
        ---Purpose: Defines the "map from" and the "map to" of the drawer.
        --          The "map from" is defined by the viewmapping.
        --          The "map to" is defined by the device.
        --          example : the X window for a X driver.

        Values (me; XF, YF, SF, XT, YT, ST, ZF: out ShortReal from Standard)
                is static;
        ---Level: Internal
        ---Purpose: Returns the "map from" and the "map to".

        --------------------------------------------
        -- Category: Methods to manage the highlight
        --------------------------------------------

        SetOverride (me: mutable; aValue: Boolean from Standard)
                is static;
        ---Level: Internal
        ---Purpose: Manages the highlight, if the highlight color index
        --          is defined (No default value)
        ---Category: Methods to manage the highlight

        SetOverrideColor (me: mutable; anIndex: Integer from Standard)
                is static;
        ---Level: Internal
        ---Purpose: Sets the highlight color index.
        --  Warning: No default value.
        ---Category: Methods to manage the highlight

        SetOffSet (me: mutable;
                anOffSet: Integer from Standard)
                is static;
        ---Level: Internal
        ---Purpose: Specifies an offset applied to the original color
        --      index when drawing a primitives, those already created
        --      and the future one.
        --  Warning: To reset the real color of the primitives when drawing
        --      then this method is called with <anOffSet> = 0.

        ---------------------------------------------
        -- Category: Methods to manage the attributes
        ---------------------------------------------

        SetLineAttrib (me: mutable;
                ColorIndex: Integer from Standard;
                TypeIndex: Integer from Standard;
                WidthIndex: Integer from Standard)
        ---Level: Internal
        ---Purpose: Methods to define the Current Line Attributes
        --  Warning: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is virtual;

        SetMarkerAttrib (me: mutable;
                ColorIndex: Integer from Standard;
                WidthIndex: Integer from Standard;
                FillMarker: Boolean from Standard)
        ---Level: Internal
        ---Purpose: Methods to define the Current Marker Attributes
        --  Warning: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;

        SetPolyAttrib (me: mutable;
                ColorIndex: Integer from Standard;
                TileIndex: Integer from Standard;
                DrawEdge: Boolean from Standard)
        ---Level: Internal
        ---Purpose: Methods to define the Current polygon Attributes
        --  Warning: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;

        SetHidingPolyAttrib (me: mutable;
                HidingColorIndex: Integer from Standard;
                FrameColorIndex: Integer from Standard;
                FrameTypeIndex: Integer from Standard;
                FrameWidthIndex: Integer from Standard)
        ---Level: Internal
        ---Purpose: Methods to define the Current hiding polygon Attributes
        --  Warning: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;

        SetTextAttrib (me: mutable;
                ColorIndex: Integer from Standard;
                FontIndex: Integer from Standard;
                aSlant: ShortReal from Standard;
                aHScale,aWScale: ShortReal from Standard;
                isUnderlined: Boolean from Standard)
        ---Level: Internal
        ---Purpose: Methods to define the Current Text Attributes
        --  Warning: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
 
        SetHidingTextAttrib (me: mutable;
                ColorIndex: Integer from Standard;
                HidingColorIndex: Integer from Standard;
                FrameColorIndex: Integer from Standard;
                FrameWidthIndex: Integer from Standard;
                FontIndex: Integer from Standard;
                aSlant: ShortReal from Standard;
                aHScale,aWScale: ShortReal from Standard;
                isUnderlined: Boolean from Standard)
        ---Level: Internal
        ---Purpose: Methods to define the Current Hiding Text Attributes
        --  Warning: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
 
        SetFramedTextAttrib (me: mutable;
                ColorIndex: Integer from Standard;
                FrameColorIndex: Integer from Standard;
                FrameWidthIndex: Integer from Standard;
                FontIndex: Integer from Standard;
                aSlant: ShortReal from Standard;
                aHScale,aWScale: ShortReal from Standard;
                isUnderlined: Boolean from Standard)
        ---Level: Internal
        ---Purpose: Methods to define the Current Framed Text Attributes
        --  Category: Methods to manage the attributes
        --  Warning: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;

        -----------------------------------------
        -- Category: Methods to manage the images
        -----------------------------------------

        IsKnownImage (me: mutable; anImageId: Transient from Standard)
        returns Boolean from Standard
        ---Level: Internal
        ---Purpose: Returns Standard_True if the associated driver
        --          have stored the image and Standard_False if not.
        --          For example, returns Standard_True if the associated
        --          driver is a X Driver.
        --  Category: Methods to manage the images
        --  Warning: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;

        ClearImage (me: mutable; anImageId: Transient from Standard)
        ---Level: Internal
        ---Purpose: Clears the image in the associated driver.
        --  Category: Methods to manage the images
        --  Warning: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;

        DrawImage (me: mutable; anImageId: Transient from Standard;
                aX, aY: ShortReal from Standard)
        ---Level: Internal
        ---Purpose: Draws the image in the associated driver.
        --          <aX>, <aY> is the center of the image.
        --  Category: Methods to manage the images
        --  Warning: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;

        ClearImageFile (me: mutable; aName: CString from Standard)
        ---Level: Internal
        ---Purpose: Clears the image file in the associated driver.
        --  Category: Methods to manage the images
        --  Warning: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;

        DrawImageFile (me: mutable; aName: CString from Standard;
                aX, aY: ShortReal from Standard;
                aScale: Factor from Quantity)
        ---Level: Internal
        ---Purpose: Draws the image in the associated driver.
        --          <aX>, <aY> is the center of the image.
        --          <aScale> = (if the image is zoomable)
        --              initial scale factor of the image *
        --              scale factor of the view.
        --          <aScale> = (if the image is not zoomable)
        --              initial scale factor of the image
        --  Category: Methods to manage the images
        --  Warning: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;

        FillAndDrawImage (me: mutable; anImageId: Transient from Standard;
                aX, aY: ShortReal from Standard;
                aWidth, aHeight: Integer from Standard;
                anArrayOfPixels: Address from Standard)
        ---Level: Internal
        ---Purpose: Stores a complete image and draws it in the associated
        --          driver.
        --          <aX>, <aY> is ????
        --  Category: Methods to manage the images
        --  Warning: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;

        FillAndDrawImage (me: mutable; anImageId: Transient from Standard;
                aX, aY: ShortReal from Standard;
                anIndexOfLine, aWidth, aHeight: Integer from Standard;
                anArrayOfPixels: Address from Standard)
        ---Level: Internal
        ---Purpose: Stores a line of an image and draws it in the associated
        --          driver.
        --          <aX>, <aY> is ????
        --  Category: Methods to manage the images
        --  Warning: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;

        ----------------------------
        -- Category: Convert methods
        ----------------------------

        GetMapFrom (me; x1, y1: ShortReal from Standard;
                x2, y2: out ShortReal from Standard)
                is static;
        ---Level: Internal
        ---Purpose: 
        --  Category: Convert methods

        GetMapFromTo (me; x1, y1: ShortReal from Standard;
                x2, y2: out ShortReal from Standard)
                is static;
        ---Level: Internal
        ---Purpose: 
        ---Category: Convert methods

        GetTextSize (me; aText: ExtendedString from TCollection;
                         aWidth,aHeight: out ShortReal from Standard)
                returns Boolean from Standard is virtual;
        ---Level: Internal
        ---Purpose: Get text size in world space with the current text
        --         attributes and returns TRUE if the driver is enabled 
        --         to get the right size (WindowDriver ONLY!). 
        --  Category: Convert methods

        GetTextSize (me; aText: ExtendedString from TCollection;
                         aWidth,aHeight,anXoffset,anYoffset: out ShortReal from Standard)
                returns Boolean from Standard is static;
        ---Level: Internal
        ---Purpose: Get text size and offsets 
        --         in world space with the current text
        --         attributes and returns TRUE if the driver is enabled 
        --         to get the right size (WindowDriver ONLY!). 
        --          NOTE that the text offsets defines the relative position of the
        --         of the text string origin from the lower left corner of the text
        --         boundary limits.
        --  Warning : SetTextAttrib(...) must be call before.
        --  Category: Convert methods

        GetFontSize (me; aHeight,aBheight,aSlant: out ShortReal from Standard)
                returns Boolean from Standard is static;
        ---Level: Internal
        ---Purpose: Get font height,baseline height and slant
        --         in world space with the current text
        --         attributes and returns TRUE if the driver is enabled 
        --       to get the right size (WindowDriver ONLY!). 
        --  Warning : SetTextAttrib(...) must be call before.
        --  Category: Convert methods

        GetImageSize (me; aFileName: CString from Standard;
                         aWidth,aHeight: out ShortReal from Standard)
                returns Boolean from Standard is static;
        ---Level: Internal
        ---Purpose: Get image size in world space 
        --         and returns TRUE if the driver is enabled 
        --         to get the right size (WindowDriver ONLY!). 
        ---Category: Convert methods

        GetImageSize (me; aFileName: CString from Standard;
                         aWidth,aHeight: out Integer from Standard)
                returns Boolean from Standard is static;
        ---Level: Internal
        ---Purpose: Get image size in pixel space 
        --         and returns TRUE if the driver is enabled 
        --         to get the right size (WindowDriver ONLY!). 
        ---Category: Convert methods

        UnMapFromTo (me;
                x1, y1: ShortReal from Standard;
                x2, y2: out ShortReal from Standard)
                is static;
        ---Level: Internal
        ---Purpose: 
        ---Category: Convert methods

        Convert (me; aValue: ShortReal from Standard)
                returns ShortReal from Standard
                is static;
        ---Level: Internal
        ---Purpose: 
        ---Category: Convert methods

        Convert (me; aValue: Integer from Standard)
                returns ShortReal from Standard
                is static;
        ---Level: Internal
        ---Purpose: 
        ---Category: Convert methods

        ConvertMapToFrom (me; x: ShortReal from Standard)
                returns ShortReal from Standard
                is static;
        ---Level: Internal
        ---Purpose: 
        ---Category: Convert methods

        Scale (me)
                returns ShortReal from Standard
                is static;
        ---Level: Internal
        ---Purpose: 
        ---Category: Convert methods

        -------------------------
        -- Category: Draw methods
        -------------------------

        DrawSegment (me : mutable; 
                x1, y1, x2, y2: ShortReal from Standard)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Level: Internal
        ---Category: Draw methods

        DrawPolyline (me : mutable;
                aDeltaX, aDeltaY: Real from Standard;
                aListX, aListY: Array1OfShortReal from TShort)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Level: Internal
        ---Category: Draw methods

        DrawPolygon (me : mutable;
                aDeltaX, aDeltaY: Real from Standard;
                aListX, aListY: Array1OfShortReal from TShort)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Level: Internal 
        ---Category: Draw methods

        DrawArc (me : mutable; 
                aDeltaX, aDeltaY: Real from Standard;
                aRadius, angle1, angle2: ShortReal from Standard)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Level: Internal
        ---Category: Draw methods
 
        DrawPolyArc (me : mutable; 
                aDeltaX, aDeltaY: Real from Standard;
                aRadius, angle1, angle2: ShortReal from Standard)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Level: Internal
        ---Category: Draw methods

        DrawInfiniteLine (me : mutable; 
                x, y, dx, dy: ShortReal from Standard)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Level: Internal
        ---Category: Draw methods

        DrawMarker (me : mutable;
                anindex: Integer from Standard;
                x, y, awidth, anheight, angle: ShortReal from Standard)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Level: Internal
        ---Category: Draw methods

        DrawText (me : mutable; 
                aText: ExtendedString from TCollection;
                x, y, angle : ShortReal from Standard;
                aType: TypeOfText from Aspect)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Level: Internal
        ---Category: Draw methods

        DrawPolyText (me : mutable; 
                aText: ExtendedString from TCollection;
                x, y, angle, margin : ShortReal from Standard;
                aType: TypeOfText from Aspect)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Level: Internal
        ---Category: Draw methods

        DrawFramedText (me : mutable; 
                aText: ExtendedString from TCollection;
                x, y, angle, margin : ShortReal from Standard;
                aType: TypeOfText from Aspect)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Level: Internal
        ---Category: Draw methods

        -------------------------------------------
        -- Category: Convert methods for primitives
        -------------------------------------------

        MapInfiniteLineFromTo (me : mutable;
                 x, y, dx, dy: ShortReal from Standard)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Level: Internal
        ---Category: Convert methods for primitives

        MapSegmentFromTo (me : mutable; 
                x1, y1, x2, y2: ShortReal from Standard;
                                aMode: Integer from Standard = 0)
        ---Level: Internal
        ---Purpose:  RRaises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is virtual;
        ---Category: Convert methods for primitives

        MapMarkerFromTo (me : mutable;
                anindex: Integer from Standard;
                x, y, awidth, anheight, angle: ShortReal from Standard;
                                aMode: Integer from Standard = 0)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Level: Internal
        ---Category: Convert methods for primitives
    	
        MapMarkersFromTo (me : mutable;
                    	 index: Integer from Standard;
                         x, y : HArray1OfShortReal from TShort;
                         awidth, anheight, angle: ShortReal from Standard;
                         aMode: Integer from Standard = 0)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Level: Internal
        ---Category: Convert methods for primitives


        MapPolylineFromTo (me : mutable;
                aListX, aListY: Array1OfShortReal from TShort;
                aNumber: Integer from Standard = 0)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Level: Internal
        ---Category: Convert methods for primitives

        MapPolylineFromTo (me : mutable; 
                x, y: ShortReal from Standard;
                aMode: Integer from Standard = 0)
        ---Level: Internal
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Category: Convert methods for primitives

        MapPolygonFromTo (me : mutable;
                aListX, aListY: Array1OfShortReal from TShort;
                aNumber: Integer from Standard = 0)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Level: Internal
        ---Category: Convert methods for primitives

        MapPolygonFromTo (me : mutable; 
                x, y: ShortReal from Standard;
                aMode: Integer from Standard = 0)
        ---Level: Internal
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Category: Convert methods for primitives

        MapTextFromTo (me : mutable; 
                aText: ExtendedString from TCollection;
                x, y, angle, aDeltax, aDeltay: ShortReal from Standard;
                aType: TypeOfText from Aspect)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is virtual;
        ---Level: Internal
        ---Category: Convert methods for primitives

        MapPolyTextFromTo (me : mutable; 
                aText: ExtendedString from TCollection;
                x, y, angle, margin, aDeltax, aDeltay: ShortReal from Standard;
                aType: TypeOfText from Aspect)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Level: Internal
        ---Category: Convert methods for primitives

        MapFramedTextFromTo (me : mutable; 
                aText: ExtendedString from TCollection;
                x, y, angle, margin, aDeltax, aDeltay: ShortReal from Standard;
                aType: TypeOfText from Aspect)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Level: Internal
        ---Category: Convert methods for primitives

        MapArcFromTo (me : mutable;
                x, y, aRadius, angle1, angle2: ShortReal from Standard;
                                aMode: Integer from Standard = 0)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is virtual;
        ---Level: Internal
        ---Category: Convert methods for primitives

        MapPolyArcFromTo (me : mutable;
                x, y, aRadius, angle1, angle2: ShortReal from Standard;
                                aMode: Integer from Standard = 0)
        ---Purpose: Raises DrawerDefinitionError if the
        --          associated driver is not defined.
        raises DrawerDefinitionError from Graphic2d is static;
        ---Level: Internal
        ---Category: Convert methods for primitives

        -----------------------------
        -- Category: Rejection method
        -----------------------------

        SetRejection (me : mutable; aClipFlag: Boolean from Standard) is static;
        ---Level: Internal
        ---Purpose: Sets the clipping flag with <aClipFlag> value.

        IsIn (me; aMinX, aMaxX, aMinY, aMaxY: ShortReal from Standard)
                returns Boolean from Standard
                is static;
        ---Level: Internal
        ---Purpose: Returns Standard_True if the given min max intersects
        --          with the drawer space.
        --          Called by the method Draw of a primitive.
        --          IsIn permits the rejection of the primitive only
        --          if the Clipping flag is TRUE.
        --          When the Clipping flag is FALSE,this method returns
        --          always TRUE.
        ---Category: Rejection method

fields
        myXF:   ShortReal from Standard;
        myYF:   ShortReal from Standard;
        mySF:   ShortReal from Standard;

        myXT:   ShortReal from Standard;
        myYT:   ShortReal from Standard;
        myST:   ShortReal from Standard;
        myZF:   ShortReal from Standard;

        myDrawPrecision:                ShortReal from Standard is protected;
        myDeflectionCoefficient:        Real from Standard is protected;
        myTypeOfDeflection:             TypeOfDeflection from Aspect is protected;
        myTextPrecision:                ShortReal from Standard;

        myOverrideColor:        Integer from Standard;
        myOverride:             Boolean from Standard;

        myOffSet:               Integer from Standard;

        -- Space of the drawing area;
        mySpaceWidth:           ShortReal from Standard is protected;
        mySpaceHeight:          ShortReal from Standard is protected;

        myDriver:               DriverPtr from Aspect is protected;
        myDriverIsDefined:      Boolean from Standard is protected;
        myWDriver:              WindowDriverPtr from Aspect is protected;
        myPDriver:              PlotterDriverPtr from PlotMgt is protected;
        myMinMaxIsActivated:    Boolean from Standard is protected;
        myMinX,myMinY,myMaxX,myMaxY : ShortReal from Standard is protected;
        myClippingIsActivated:    Boolean from Standard is protected;

end Drawer from Graphic2d;

