-- File:        PersonAndOrganization.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWPersonAndOrganization from RWStepBasic

	---Purpose : Read & Write Module for PersonAndOrganization

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     PersonAndOrganization from StepBasic,
     EntityIterator from Interface

is

	Create returns RWPersonAndOrganization;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable PersonAndOrganization from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : PersonAndOrganization from StepBasic);

	Share(me; ent : PersonAndOrganization from StepBasic; iter : in out EntityIterator);

end RWPersonAndOrganization;
