-- File:	TopoDS_Edge.cdl
-- Created:	Mon Dec 17 10:48:25 1990
-- Author:	Remi Lequette
---Copyright:	 Matra Datavision 1990, 1992


class Edge from TopoDS inherits Shape

	---Purpose: Describes an edge which
-- - references an underlying edge with the potential to
--   be given a location and an orientation
-- - has a location for the underlying edge, giving its
--   placement in the local coordinate system
-- - has an orientation for the underlying edge, in terms
--   of its geometry (as opposed to orientation in
--   relation to other shapes).

is
    Create returns Edge from TopoDS;
    ---C++: inline
	---Purpose: Undefined Edge.

end Edge;
