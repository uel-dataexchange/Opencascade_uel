-- File:	GCPnts_QuasiUniformDeflection.cdl
-- Created:	Thu Nov  2 14:57:07 1995
-- Author:	Jacques GOUSSARD
--		<jag@bravox>
---Copyright:	 Matra Datavision 1995


class QuasiUniformDeflection from GCPnts 

    ---Purpose: This  class computes  a  distribution of  points  on a
    --          curve. The points may respect the deflection. The algorithm
    --          is not based on the  classical prediction (with second
    --          derivative of curve), but either  on the evaluation of
    --          the distance between the   mid point and the  point of
    --          mid parameter of    the two points,   or  the distance
    --          between the mid point and  the point at parameter  0.5
    --          on the cubic interpolation of the two points and their
    --          tangents.
    -- Note: this algorithm is faster than a
    -- GCPnts_UniformDeflection algorithm, and is
    -- able to work with non-"C2" continuous curves.
    -- However, it generates more points in the distribution.
        
uses 
    Pnt            from gp,
    Curve          from Adaptor3d,
    Curve2d        from Adaptor2d,
    Shape          from GeomAbs,
    SequenceOfPnt  from TColgp,
    SequenceOfReal from TColStd
    

raises DomainError       from Standard, 
       ConstructionError from Standard,
       OutOfRange        from Standard,
       NotDone           from StdFail

is
        
    Create 
    	---Purpose: Constructs an empty algorithm. To define the problem
        -- to be solved, use the function Initialize.
    	returns QuasiUniformDeflection from GCPnts;

    Create(C : in out Curve from Adaptor3d; Deflection : Real; 
           Continuity: Shape  from  GeomAbs  =  GeomAbs_C1)
        --- Purpose : Computes  a QuasiUniform Deflection distribution
        --  of points on the Curve <C>.
    	returns QuasiUniformDeflection from GCPnts
     	raises ConstructionError;

    Create(C : in out Curve2d from Adaptor2d; Deflection : Real; 
           Continuity: Shape  from  GeomAbs  =  GeomAbs_C1)
        --- Purpose : Computes  a QuasiUniform Deflection distribution
        --  of points on the Curve <C>.
    	returns QuasiUniformDeflection from GCPnts
     	raises ConstructionError;

    Create(C : in out Curve from Adaptor3d; Deflection, U1, U2 : Real; 
           Continuity: Shape  from  GeomAbs  =  GeomAbs_C1)
        --- Purpose  : Computes a QuasiUniform Deflection distribution
        --  of points on a part of the Curve <C>.
     	returns QuasiUniformDeflection from GCPnts
     	raises ConstructionError,
               DomainError;

    Create(C : in out Curve2d from Adaptor2d; Deflection, U1, U2 : Real; 
           Continuity: Shape  from  GeomAbs  =  GeomAbs_C1)
        ---Purpose :  Computes  a QuasiUniform Deflection distribution
        --  of points on a part of the Curve <C>.
	-- This and the above algorithms compute a distribution of points:
	-- -   on the curve C, or
	-- -   on the part of curve C limited by the two
	--   parameter values U1 and U2,
	-- where the deflection resulting from the distributed
	-- points is not greater than Deflection.
	-- The first point of the distribution is either the origin of
	-- curve C or the point of parameter U1. The last point
	-- of the distribution is either the end point of curve C or
	-- the point of parameter U2.
	-- Intermediate points of the distribution are built such
	-- that the deflection is not greater than Deflection.
	-- Using the following evaluation of the deflection:
	-- if Pi and Pj are two consecutive points of the
	-- distribution, respectively of parameter ui and uj on
	-- the curve, the deflection is the distance between:
	-- -   the mid-point of Pi and Pj (the center of the
	--   chord joining these two points)
	-- -   and the point of mid-parameter of these two
	--   points (the point of parameter [(ui+uj) / 2 ] on curve C).
	--   Continuity, defaulted to GeomAbs_C1, gives the
	--   degree of continuity of the curve C. (Note that C is an
	-- Adaptor3d_Curve or an Adaptor2d_Curve2d
	-- object, and does not know the degree of continuity of
	-- the underlying curve).
	-- Use the function IsDone to verify that the
	-- computation was successful, the function NbPoints
	-- to obtain the number of points of the computed
	-- distribution, and the function Parameter to read the
	-- parameter of each point.
	-- Warning
	-- -   The roles of U1 and U2 are inverted if U1 > U2.
	-- -   Derivative functions on the curve are called
	--   according to Continuity. An error may occur if
	--   Continuity is greater than the real degree of
	--   continuity of the curve.
	-- Warning
	-- C is an adapted curve, i.e. an object which is an
	-- interface between:
	-- -   the services provided by either a 2D curve from
	--   the package Geom2d (in the case of an
	--   Adaptor2d_Curve2d curve) or a 3D curve from
	--   the package Geom (in the case of an
	--   Adaptor3d_Curve curve),
	-- -   and those required on the curve by the
	--   computation algorithm.
     	returns QuasiUniformDeflection from GCPnts
     	raises ConstructionError,
               DomainError;

    Initialize(me : in out; C : in out Curve from Adaptor3d; Deflection : Real; 
           Continuity: Shape  from  GeomAbs  =  GeomAbs_C1)
    	---Purpose: Initialize the algoritms with <C>, <Deflection>
     	raises ConstructionError
	is static;

    Initialize(me : in out; C : in out Curve2d from Adaptor2d; Deflection : Real; 
           Continuity: Shape  from  GeomAbs  =  GeomAbs_C1)
    	---Purpose: Initialize the algoritms with <C>, <Deflection>
     	raises ConstructionError
	is static;

    Initialize(me : in out; C : in out Curve from Adaptor3d; Deflection, U1, U2 : Real; 
           Continuity: Shape  from  GeomAbs  =  GeomAbs_C1)
        ---Purpose: Initialize the algoritms with <C>, <Deflection>,
    	--          <U1>,<U2>
     	raises ConstructionError,
               DomainError
	is static;
  
    Initialize(me : in out; C : in out Curve2d from Adaptor2d; 
    	    	            Deflection, U1, U2 : Real; 
           Continuity: Shape  from  GeomAbs  =  GeomAbs_C1)
        ---Purpose: Initialize  the  algoritms with <C>, <Deflection>,
        --          -- <U1>,<U2>
	--    This and the above algorithms initialize (or reinitialize)
	--        this algorithm and compute a distribution of points:
	-- -   on the curve C, or
	-- -   on the part of curve C limited by the two
	--   parameter values U1 and U2,
	-- where the deflection resulting from the distributed
	-- points is not greater than Deflection.
	-- The first point of the distribution is either the origin
	-- of curve C or the point of parameter U1. The last
	-- point of the distribution is either the end point of
	-- curve C or the point of parameter U2.
	-- Intermediate points of the distribution are built in
	-- such a way that the deflection is not greater than
	-- Deflection. Using the following evaluation of the deflection:
	-- if Pi and Pj are two consecutive points of the
	-- distribution, respectively of parameter ui and uj
	-- on the curve, the deflection is the distance between:
	-- -   the mid-point of Pi and Pj (the center of the
	--   chord joining these two points)
	-- -   and the point of mid-parameter of these two
	--   points (the point of parameter [(ui+uj) / 2 ] on curve C).
	--   Continuity, defaulted to GeomAbs_C1, gives the
	-- degree of continuity of the curve C. (Note that C is
	-- an Adaptor3d_Curve or an
	-- Adaptor2d_Curve2d object, and does not know
	-- the degree of continuity of the underlying curve).
	-- Use the function IsDone to verify that the
	-- computation was successful, the function NbPoints
	-- to obtain the number of points of the computed
	-- distribution, and the function Parameter to read
	-- the parameter of each point.
	-- Warning
	-- -   The roles of U1 and U2 are inverted if U1 > U2.
	-- -   Derivative functions on the curve are called
	--   according to Continuity. An error may occur if
	--   Continuity is greater than the real degree of
	--   continuity of the curve.
	-- Warning
	-- C is an adapted curve, i.e. an object which is an
	-- interface between:
	-- -   the services provided by either a 2D curve from
	--   the package Geom2d (in the case of an
	--   Adaptor2d_Curve2d curve) or a 3D curve from
	--   the package Geom (in the case of an Adaptor3d_Curve curve),
	-- and those required on the curve by the computation algorithm.
    raises ConstructionError,
               DomainError
	is static;
  	
    IsDone(me) returns Boolean
	---C++: inline
	---	Purpose:
	-- Returns true if the computation was successful.
	-- IsDone is a protection against:
	-- -   non-convergence of the algorithm
	-- -   querying the results before computation.
    	is static;
	       
    NbPoints(me) returns Integer
	---C++: inline
	---Purpose:
	-- Returns the number of points of the distribution
	-- computed by this algorithm.
	-- Exceptions
	-- StdFail_NotDone if this algorithm has not been
	-- initialized, or if the computation was not successful.
    	is static;
  
    Parameter(me; Index : Integer) returns Real 
	---C++: inline
        --- Purpose : Returns the parameter of the point of index Index in
	-- the distribution computed by this algorithm.
	-- Warning
	-- Index must be greater than or equal to 1, and less
	-- than or equal to the number of points of the
	-- distribution. However, pay particular attention as this
	-- condition is not checked by this function.
	-- Exceptions
	-- StdFail_NotDone if this algorithm has not been
	-- initialized, or if the computation was not successful.
    	is static;
	
    Value(me; Index : Integer) returns Pnt from gp 
        --- Purpose : Returns the point of index Index in the distribution
	-- computed by this algorithm.
	-- Warning
	-- Index must be greater than or equal to 1, and less
	-- than or equal to the number of points of the
	-- distribution. However, pay particular attention as this
	-- condition is not checked by this function.
	-- Exceptions
	-- StdFail_NotDone if this algorithm has not been
	-- initialized, or if the computation was not successful.
    	is static;
    
    Deflection(me) returns Real
	---C++: inline
      	--- Purpose : Returns the deflection between the curve and the
	-- polygon resulting from the points of the distribution
	-- computed by this algorithm.
	-- This is the value given to the algorithm at the time
	-- of construction (or initialization).
	-- Exceptions
	-- StdFail_NotDone if this algorithm has not been
	-- initialized, or if the computation was not successful.
	is static;

fields

    myDone          : Boolean;
    myDeflection    : Real;
    myParams        : SequenceOfReal from TColStd;
    myPoints        : SequenceOfPnt  from TColgp;
    myCont          : Shape          from GeomAbs;
    
end QuasiUniformDeflection;

