-- File:        LoopAndPath.cdl
-- Created:     Mon Dec  4 12:02:37 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWLoopAndPath from RWStepShape

	---Purpose : Read & Write Module for LoopAndPath

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     LoopAndPath from StepShape,
     EntityIterator from Interface

is

	Create returns RWLoopAndPath;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable LoopAndPath from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : LoopAndPath from StepShape);

	Share(me; ent : LoopAndPath from StepShape; iter : in out EntityIterator);

end RWLoopAndPath;
