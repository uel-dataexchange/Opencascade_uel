-- File:	RWStepBasic_RWContractAssignment.cdl
-- Created:	Fri Nov 26 16:26:37 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWContractAssignment from RWStepBasic

    ---Purpose: Read & Write tool for ContractAssignment

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ContractAssignment from StepBasic

is
    Create returns RWContractAssignment from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ContractAssignment from StepBasic);
	---Purpose: Reads ContractAssignment

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ContractAssignment from StepBasic);
	---Purpose: Writes ContractAssignment

    Share (me; ent : ContractAssignment from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWContractAssignment;
