-- File:	MakeArcOfParabola.cdl
-- Created:	Mon Sep 28 11:51:03 1992
-- Author:	Remi GILET
--		<reg@sdsun2>
---Copyright:	 Matra Datavision 1992

class MakeArcOfParabola from GCE2d inherits Root from GCE2d
    	---Purpose: Implements construction algorithms for an arc of
    	-- parabola in the plane. The result is a Geom2d_TrimmedCurve curve.
    	-- A MakeArcOfParabola object provides a framework for:
    	-- -   defining the construction of the arc of parabola,
    	-- -   implementing the construction algorithm, and
    	-- -   consulting the results. In particular, the Value
    	--   function returns the constructed arc of parabola.
        
uses Pnt2d        from gp,
     Parab2d      from gp,
     Real         from Standard,
     Boolean      from Standard,
     TrimmedCurve from Geom2d

raises NotDone from StdFail

is

Create(Parab          : Parab2d from gp                      ;
       Alpha1, Alpha2 : Real    from Standard                ;
       Sense          : Boolean from Standard = Standard_True) 
    returns MakeArcOfParabola;
    	---Purpose: Make an arc of Parabola (TrimmedCurve from Geom2d) from 
    	--          a Parabola between two parameters Alpha1 and Alpha2.

Create(Parab : Parab2d from gp                      ;
       P     : Pnt2d   from gp                      ;
       Alpha : Real    from Standard                ;
       Sense : Boolean from Standard = Standard_True)
    returns MakeArcOfParabola;
    	---Purpose: Make an arc of Parabola (TrimmedCurve from Geom2d) from 
    	--          a Parabola between point <P> and the parameter
        --          Alpha.

Create(Parab : Parab2d from gp                      ;
       P1    : Pnt2d   from gp                      ;
       P2    : Pnt2d   from gp                      ;
       Sense : Boolean from Standard = Standard_True) 
    returns MakeArcOfParabola;
    	---Purpose: Make an arc of Parabola (TrimmedCurve from Geom2d) from 
    	--          a Parabola between two points P1 and P2.
    	-- Please, note: the orientation of the arc of parabola is:
    	--   -   the trigonometric sense if Sense is not defined
    	--    or is true (default value), or
    	--   -   the opposite sense if Sense is false.
    	-- - IsDone always returns true.
        
Value(me) returns TrimmedCurve from Geom2d
    raises NotDone
    is static;
    	---C++: return const&
    	---Purpose: Returns the constructed arc of parabola.
    
Operator(me) returns TrimmedCurve from Geom2d
    is static;
    	---C++: return const&
    	---C++: alias "Standard_EXPORT operator Handle_Geom2d_TrimmedCurve() const;"

fields

    TheArc : TrimmedCurve from Geom2d;
    --The solution from Geom2d.
    
end MakeArcOfParabola;
