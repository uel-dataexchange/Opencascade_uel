-- File:	IGESGeom_ToolBoundary.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolBoundary  from IGESGeom

    ---Purpose : Tool to work on a Boundary. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses Boundary from IGESGeom,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolBoundary;
    ---Purpose : Returns a ToolBoundary, ready to work


    ReadOwnParams (me; ent : mutable Boundary;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : Boundary;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : Boundary;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a Boundary <ent>, from
    --           its specific (own) parameters

    OwnCorrect (me; ent : mutable Boundary) returns Boolean  is static;
    ---Purpose : Sets automatic unambiguous Correction on a Boundary
    --           (if BoundaryType = 0, Nullify all ParameterCurves)

    DirChecker (me; ent : Boundary) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : Boundary;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : Boundary; entto : mutable Boundary;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : Boundary;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolBoundary;
