-- File:	Geom2dAPI.cdl
-- Created:	Wed Mar 23 15:00:46 1994
-- Author:	Bruno DUMORTIER
--		<dub@fuegox>
---Copyright:	 Matra Datavision 1994

package Geom2dAPI

	---Purpose: The  Geom2dAPI  package  provides  an  Application
	--          Programming Interface for the Geometry.
	--          
	--          The API is a set of classes aiming to provide :
	--          
	--          * High level and simple calls  for the most common
	--          operations. 
	--          
	--          *    Keeping   an   access  on    the    low-level
	--          implementation of high-level calls.
	--          
	-- 	    
	-- 	    The API  provides classes to  call the algorithmes
	-- 	    of the Geometry
	-- 	    
	-- 	    * The  constructors  of the classes  provides  the
	-- 	    different constructions methods.
	-- 	    
	-- 	    * The  class keeps as fields the   different tools
	-- 	    used by the algorithmes
	-- 	    
	-- 	    *   The class  provides  a  casting  method to get
	-- 	    automatically the  result  with  a   function-like
	-- 	    call. 
	-- 	    
	-- 	    For example to evaluate the distance <D> between a
	-- 	    point <P> and a curve <C>, one can writes :
	-- 	    
	-- 	        D = Geom2dAPI_ProjectPointOnCurve(P,C);
	-- 	    
	-- 	    or
	-- 	    
	-- 	        Geom2dAPI_ProjectPointOnCurve PonC(P,C);
	-- 	        D = PonC.LowerDistance();
	-- 	    


uses

    Geom2d,
    gp,
    TColgp,
    Extrema,
    Geom2dAdaptor,
    Geom2dInt,
    GeomAbs,
    TColStd,
    Quantity, 
    Approx,
    StdFail
    

is

    ------------------------------------------------------------------
    -- This classes  provides algo  to  evaluate  the distance between
    -- points and curves, curves and curves. 
    ------------------------------------------------------------------

    class ProjectPointOnCurve;

    class ExtremaCurveCurve;
    


    ------------------------------------------------------------------
    -- This classes provides algo to evaluate a curve  passing through
    -- an array of points.
    ------------------------------------------------------------------

    --- Approximation:
    --  
    class PointsToBSpline;
    
    
    --- Interpolation:
    --
    class Interpolate;
    
    
    ------------------------------------------------------------------
    -- This classes provides algo to evaluate an intersection between 
    -- two 2d-Curves.
    ------------------------------------------------------------------

    class InterCurveCurve;


end Geom2dAPI;
