-- File:	BRepOffsetAPI_MakeOffset.cdl
-- Created:	Mon Sep 18 13:40:56 1995
-- Author:	Bruno DUMORTIER
--		<dub@fuegox>
---Copyright:	 Matra Datavision 1995


class MakeOffset from BRepOffsetAPI inherits MakeShape from BRepBuilderAPI

	---Purpose: Describes algorithms for offsetting wires from a set of
    	-- wires contained in a planar face.
    	-- A MakeOffset object provides a framework for:
    	-- - defining the construction of an offset,
    	-- - implementing the construction algorithm, and
    	-- - consulting the result. 

uses
    Shape             from TopoDS,
    Wire              from TopoDS,
    Face              from TopoDS,
    ListOfShape       from TopTools,
    OffsetWire        from BRepFill, 
    ListOfOffsetWire  from BRepFill,
    JoinType          from GeomAbs
    
    
raises
    ConstructionError from Standard
    
is
    Create returns MakeOffset from BRepOffsetAPI;
    	---Purpose: Constructs an algorithm for creating an empty offset
    Create( Spine : Face from TopoDS;
    	    Join  : JoinType from GeomAbs = GeomAbs_Arc)
    returns MakeOffset from BRepOffsetAPI;
    	---Purpose: Constructs an algorithm for creating an algorithm
    	-- to build parallels to the spine Spine   
    Init( me    : in out;
    	  Spine : Face     from TopoDS; 
    	  Join  : JoinType from GeomAbs  =  GeomAbs_Arc)
	---Purpose: Initializes the algorithm to construct parallels to the spine Spine.
    	-- Join defines the type of parallel generated by the
    	-- salient vertices of the spine. The default type is
    	-- GeomAbs_Arc where the vertices generate sections
    	-- of a circle. At present, this is the only construction type implemented.
    is static;
    
    Create( Spine : Wire from TopoDS;
    	    Join  : JoinType from GeomAbs = GeomAbs_Arc)
    returns MakeOffset from BRepOffsetAPI;
    
    Init( me    : in out;
    	  Join  : JoinType from GeomAbs  =  GeomAbs_Arc)
	---Purpose: Initialize the evaluation of Offseting.
    is static;

    AddWire (me : in out;
    	     Spine : Wire from TopoDS)
        ---Purpose: Initializes the algorithm to construct parallels to the wire Spine.
    is static;

    Perform (me : in out; 
    	     Offset : Real from Standard;
    	     Alt    : Real from Standard = 0.0)
	---Purpose:  Computes a parallel to the spine at distance Offset and
    	-- at an altitude Alt from the plane of the spine in relation
    	-- to the normal to the spine.
    	-- Exceptions: Standard_ConstructionError if the offset is not built.
    raises
    	ConstructionError from Standard
    is static;

	
    Build(me : in out)
    is redefined;
	---Purpose: Builds the resulting shape (redefined from MakeShape).
	---Level: Public    

    Generated  (me: in out; S : Shape from TopoDS)
    	---Purpose: returns a list of the created shapes
    	--          from the shape <S>.
    	---C++:     return const &
	---Level: Public
    returns ListOfShape from TopTools
    is redefined;


fields

    myIsInitialized : Boolean          from Standard;
    myLastIsLeft    : Boolean          from Standard;
    myJoin          : JoinType         from GeomAbs;	
    myFace          : Face             from TopoDS;
    myWires         : ListOfShape      from TopTools;   
    myLeft          : ListOfOffsetWire from BRepFill;
    myRight         : ListOfOffsetWire from BRepFill;
    
end MakeOffset;
