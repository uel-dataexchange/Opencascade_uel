-- File:	RWStepShape_RWDimensionalSizeWithPath.cdl
-- Created:	Tue Apr 18 16:42:58 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWDimensionalSizeWithPath from RWStepShape

    ---Purpose: Read & Write tool for DimensionalSizeWithPath

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    DimensionalSizeWithPath from StepShape

is
    Create returns RWDimensionalSizeWithPath from RWStepShape;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : DimensionalSizeWithPath from StepShape);
	---Purpose: Reads DimensionalSizeWithPath

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: DimensionalSizeWithPath from StepShape);
	---Purpose: Writes DimensionalSizeWithPath

    Share (me; ent : DimensionalSizeWithPath from StepShape;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWDimensionalSizeWithPath;
