-- File:	RWStepFEA_RWFeaCurveSectionGeometricRelationship.cdl
-- Created:	Wed Jan 22 17:31:43 2003 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFeaCurveSectionGeometricRelationship from RWStepFEA

    ---Purpose: Read & Write tool for FeaCurveSectionGeometricRelationship

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FeaCurveSectionGeometricRelationship from StepFEA

is
    Create returns RWFeaCurveSectionGeometricRelationship from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FeaCurveSectionGeometricRelationship from StepFEA);
	---Purpose: Reads FeaCurveSectionGeometricRelationship

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FeaCurveSectionGeometricRelationship from StepFEA);
	---Purpose: Writes FeaCurveSectionGeometricRelationship

    Share (me; ent : FeaCurveSectionGeometricRelationship from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFeaCurveSectionGeometricRelationship;
