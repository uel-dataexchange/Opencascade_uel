-- File:	RWStepFEA_RWFeaMaterialPropertyRepresentation.cdl
-- Created:	Thu Dec 12 17:51:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFeaMaterialPropertyRepresentation from RWStepFEA

    ---Purpose: Read & Write tool for FeaMaterialPropertyRepresentation

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FeaMaterialPropertyRepresentation from StepFEA

is
    Create returns RWFeaMaterialPropertyRepresentation from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FeaMaterialPropertyRepresentation from StepFEA);
	---Purpose: Reads FeaMaterialPropertyRepresentation

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FeaMaterialPropertyRepresentation from StepFEA);
	---Purpose: Writes FeaMaterialPropertyRepresentation

    Share (me; ent : FeaMaterialPropertyRepresentation from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFeaMaterialPropertyRepresentation;
