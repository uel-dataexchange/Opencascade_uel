-- File:	Prs3d_Line.cdl
-- Created:	Wed Dec 16 12:39:30 1992
-- Author:	Jean Louis FRENKEL
--		<jlf@mastox>
---Copyright:	 Matra Datavision 1992

generic class Line from Prs3d 
                            (anyLine as any; 
    	    	    	     LineTool as any) -- as LineTool from Prs3d
inherits Root from Prs3d

---Purpose: draws a broken line.
--          
          
uses 
    Presentation from Prs3d,
    Drawer from Prs3d,
    TypeOfLinePicking from Prs3d,
    Length from Quantity
    
is
    Add(myclass; aPresentation: Presentation from Prs3d; 
         	 aLine: anyLine;
    	    	 aDrawer: Drawer from Prs3d);
		 
    ---Purpose: adds to the presentation aPresentation the drawing of the
    --          broken line aLine.     
    --          The aspect is defined by LineAspect in aDrawer.


    Add(myclass; aPresentation: Presentation from Prs3d; 
         	 aLine: anyLine);
    
    ---Purpose: adds to the presentation aPresentation the drawing of the
    --          broken line aLine.     
    --          The aspect is the current aspect.



    Pick(myclass; X,Y,Z: Length from Quantity;
    	          aDistance: Length from Quantity;
                  aLine: anyLine;
    	          aDrawer: Drawer from Prs3d;
                  TypeOfPicking: TypeOfLinePicking from Prs3d)
    returns Integer from Standard;

    ---Purpose: if TypeOfLinePicking is set to Prs3d_TOLP_Point
    --          returns the number of the point the most near of the 
    --          point (X,Y,Z). The distance between the point and
    --          (X,Y,Z) must be less then aDistance. If no point corresponds,
    --          0 is returned.
    --          if TypeOfLinePicking is set to Prs3d_TOLP_Segment returns
    --          the number of the segment the most near of the point (X,Y,Z).
    --          The distance between the segment and (X,Y,Z) must be less 
    --          then aDistance. If no segment corresponds, 0 is returned.


end Line;
