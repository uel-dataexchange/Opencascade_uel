-- File:        Axis1Placement.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWAxis1Placement from RWStepGeom

	---Purpose : Read & Write Module for Axis1Placement

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     Axis1Placement from StepGeom,
     EntityIterator from Interface

is

	Create returns RWAxis1Placement;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable Axis1Placement from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : Axis1Placement from StepGeom);

	Share(me; ent : Axis1Placement from StepGeom; iter : in out EntityIterator);

end RWAxis1Placement;
