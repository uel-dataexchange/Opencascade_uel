-- File:	IGESAppli_ToolNodalConstraint.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolNodalConstraint  from IGESAppli

    ---Purpose : Tool to work on a NodalConstraint. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses NodalConstraint from IGESAppli,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolNodalConstraint;
    ---Purpose : Returns a ToolNodalConstraint, ready to work


    ReadOwnParams (me; ent : mutable NodalConstraint;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : NodalConstraint;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : NodalConstraint;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a NodalConstraint <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : NodalConstraint) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : NodalConstraint;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : NodalConstraint; entto : mutable NodalConstraint;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : NodalConstraint;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolNodalConstraint;
