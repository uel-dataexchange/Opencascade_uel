-- File:	RWStepFEA_RWAlignedSurface3dElementCoordinateSystem.cdl
-- Created:	Thu Dec 26 15:06:35 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWAlignedSurface3dElementCoordinateSystem from RWStepFEA

    ---Purpose: Read & Write tool for AlignedSurface3dElementCoordinateSystem

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    AlignedSurface3dElementCoordinateSystem from StepFEA

is
    Create returns RWAlignedSurface3dElementCoordinateSystem from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : AlignedSurface3dElementCoordinateSystem from StepFEA);
	---Purpose: Reads AlignedSurface3dElementCoordinateSystem

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: AlignedSurface3dElementCoordinateSystem from StepFEA);
	---Purpose: Writes AlignedSurface3dElementCoordinateSystem

    Share (me; ent : AlignedSurface3dElementCoordinateSystem from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWAlignedSurface3dElementCoordinateSystem;
