-- File:        ClosedShell.cdl
-- Created:     Fri Dec  1 11:11:16 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993


class ClosedShell from StepShape 

inherits ConnectedFaceSet from StepShape 

uses

	HAsciiString from TCollection, 
	HArray1OfFace from StepShape
is

	Create returns mutable ClosedShell;
	---Purpose: Returns a ClosedShell


end ClosedShell;
