-- File:        ElementarySurface.cdl
-- Created:     Mon Dec  4 12:02:26 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWElementarySurface from RWStepGeom

	---Purpose : Read & Write Module for ElementarySurface

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ElementarySurface from StepGeom,
     EntityIterator from Interface

is

	Create returns RWElementarySurface;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ElementarySurface from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : ElementarySurface from StepGeom);

	Share(me; ent : ElementarySurface from StepGeom; iter : in out EntityIterator);

end RWElementarySurface;
