-- File:	GeomToStep_MakeElementarySurface.cdl
-- Created:	Tue Jun 22 14:24:10 1993
-- Author:	Martine LANGLOIS
--		<mla@mastox>
---Copyright:	 Matra Datavision 1993

class MakeElementarySurface from GeomToStep inherits Root from GeomToStep

    ---Purpose: This class implements the mapping between classes 
    --          ElementarySurface from Geom and the class ElementarySurface
    --          from StepGeom which describes a ElementarySurface from
    --          prostep. As ElementarySurface is an abstract Surface this
    --          class is an access to the sub-class required.
  
uses ElementarySurface from Geom,
     ElementarySurface from StepGeom
     
raises NotDone from StdFail
     
is 

Create ( S : ElementarySurface from Geom ) returns MakeElementarySurface;

Value (me) returns ElementarySurface from StepGeom
    raises NotDone
    is static;
    ---C++: return const&
 
fields

    theElementarySurface : ElementarySurface from StepGeom;
    	-- The solution from StepGeom
    	
end MakeElementarySurface;



