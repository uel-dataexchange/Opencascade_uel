-- File:	RWStepFEA_RWNodeRepresentation.cdl
-- Created:	Thu Dec 12 17:51:06 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWNodeRepresentation from RWStepFEA

    ---Purpose: Read & Write tool for NodeRepresentation

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    NodeRepresentation from StepFEA

is
    Create returns RWNodeRepresentation from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : NodeRepresentation from StepFEA);
	---Purpose: Reads NodeRepresentation

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: NodeRepresentation from StepFEA);
	---Purpose: Writes NodeRepresentation

    Share (me; ent : NodeRepresentation from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWNodeRepresentation;
