-- File:        RectangularTrimmedSurface.cdl
-- Created:     Mon Dec  4 12:02:30 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWRectangularTrimmedSurface from RWStepGeom

	---Purpose : Read & Write Module for RectangularTrimmedSurface

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     RectangularTrimmedSurface from StepGeom,
     EntityIterator from Interface

is

	Create returns RWRectangularTrimmedSurface;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable RectangularTrimmedSurface from StepGeom);

	WriteStep (me; SW : in out StepWriter; ent : RectangularTrimmedSurface from StepGeom);

	Share(me; ent : RectangularTrimmedSurface from StepGeom; iter : in out EntityIterator);

end RWRectangularTrimmedSurface;
