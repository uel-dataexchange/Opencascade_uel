-- File:	IGESGeom_ToolCompositeCurve.cdl
-- Created:	Thu Oct 14 19:16:58 1993
-- Author:	Christian CAILLET
--		<cky@bravox>
---Copyright:	 Matra Datavision 1993


class ToolCompositeCurve  from IGESGeom

    ---Purpose : Tool to work on a CompositeCurve. Called by various Modules
    --           (ReadWriteModule, GeneralModule, SpecificModule)

uses CompositeCurve from IGESGeom,
     IGESReaderData, ParamReader, IGESWriter, EntityIterator,
     DirChecker,     ShareTool,   Check,      CopyTool,   IGESDumper, Messenger from Message

raises DomainError

is

    Create returns ToolCompositeCurve;
    ---Purpose : Returns a ToolCompositeCurve, ready to work


    ReadOwnParams (me; ent : mutable CompositeCurve;
    	    	   IR : IGESReaderData; PR : in out ParamReader)
    	raises DomainError  is static;
    ---Purpose : Reads own parameters from file. <PR> gives access to them,
    --           <IR> detains parameter types and values

    WriteOwnParams (me; ent : CompositeCurve;
    	    	    IW : in out IGESWriter)  is static;
    ---Purpose : Writes own parameters to IGESWriter


    OwnShared  (me; ent : CompositeCurve;
    	        iter : in out EntityIterator)  is static;
    ---Purpose : Lists the Entities shared by a CompositeCurve <ent>, from
    --           its specific (own) parameters

    DirChecker (me; ent : CompositeCurve) returns DirChecker  is static;
    ---Purpose : Returns specific DirChecker

    OwnCheck   (me; ent : CompositeCurve;
    	        shares  : ShareTool; ach : in out Check)  is static;
    ---Purpose : Performs Specific Semantic Check


    OwnCopy    (me; entfrom : CompositeCurve; entto : mutable CompositeCurve;
    	        TC : in out CopyTool)  is static;
    ---Purpose : Copies Specific Parameters


    OwnDump (me; ent : CompositeCurve;
    	     dumper  : IGESDumper;  S : Messenger from Message; own : Integer)
        is static;
    ---Purpose : Dump of Specific Parameters

end ToolCompositeCurve;
