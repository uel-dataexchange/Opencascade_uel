-- File:        GaussMultipleIntegration.cdl
-- Created:     Tue May 14 18:22:12 1991
-- Author:      Laurent PAINNOT
--              <lpa@topsn3>
---Copyright:    Matra Datavision 1991, 1992



class GaussMultipleIntegration from math
    ---Purpose:
    -- This class implements the integration of a function of multiple 
    -- variables between the parameter bounds Lower[a..b] and Upper[a..b].
    --  Warning: Each element of Order must be inferior or equal to 61.


uses Vector from math, 
     IntegerVector from math, 
     MultipleVarFunction from math,
     OStream from Standard

raises NotDone from StdFail

is

     Create(F: in out MultipleVarFunction; Lower, Upper: Vector;
     	    Order: IntegerVector)
     ---Purpose:
     -- The Gauss-Legendre integration with Order = points of 
     -- integration for each unknow, is done on the function F 
     -- between the bounds Lower and Upper.
     
     returns GaussMultipleIntegration;
     
     IsDone(me)
     	---Purpose: returns True if all has been correctly done.
    	---C++: inline

     returns Boolean
     is static;
     
     Value(me)
     	---Purpose: returns the value of the integral.
    	---C++: inline

     returns Real
     raises NotDone
     is static;


    Dump(me; o: in out OStream)
    	---Purpose: Prints information on the current state of the object.

    is static;



fields

Val: Real;
Done: Boolean;

end GaussMultipleIntegration;
