-- File:	BinMDataXtd_ShapeDriver.cdl
-- Created:	Thu May 13 11:26:08 2004
-- Author:	Sergey ZARITCHNY <szy@opencascade.com>
-- modified     13.04.2009 Sergey Zaritchny
-- Copyright:	Open CasCade S.A. 2004

class ShapeDriver from BinMDataXtd inherits ADriver from BinMDF

        ---Purpose:  Shape attribute Driver.

uses
    MessageDriver    from CDM,
    SRelocationTable from BinObjMgt,
    RRelocationTable from BinObjMgt,
    Persistent       from BinObjMgt,
    Attribute        from TDF

is
    Create (theMessageDriver:MessageDriver from CDM)
        returns mutable ShapeDriver from BinMDataXtd;

    NewEmpty (me)  returns mutable Attribute from TDF
    	is redefined;

    Paste(me; Source     : Persistent from BinObjMgt;
              Target     : mutable Attribute from TDF;
              RelocTable : out RRelocationTable from BinObjMgt)
        returns Boolean from Standard is redefined;

    Paste(me; Source     : Attribute from TDF;
              Target     : in out Persistent from BinObjMgt;
              RelocTable : out SRelocationTable from BinObjMgt)
    	is redefined;

end ShapeDriver;

