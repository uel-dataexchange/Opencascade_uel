-- File:        MeasureWithUnit.cdl
-- Created:     Mon Dec  4 12:02:28 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWMeasureWithUnit from RWStepBasic

	---Purpose : Read & Write Module for MeasureWithUnit

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     MeasureWithUnit from StepBasic,
     EntityIterator from Interface

is

	Create returns RWMeasureWithUnit;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable MeasureWithUnit from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : MeasureWithUnit from StepBasic);

	Share(me; ent : MeasureWithUnit from StepBasic; iter : in out EntityIterator);

end RWMeasureWithUnit;
