-- File:	TestTopOpeDraw_DrawableC2D.cdl
-- Created:	Fri Dec  1 17:56:57 1995
-- Author:	Jean Yves LEBEY
--		<jyl@meteox>
---Copyright:	 Matra Datavision 1995

class DrawableC2D from TestTopOpeDraw inherits Curve2d from DrawTrSurf

uses  

    Interpretor from Draw,
    Curve from Geom2d,
    Color from Draw,
    Display from Draw,
    Text2D from Draw,
    CString from Standard,
    Pnt2d from gp

is

    Create (C : Curve from Geom2d; CColor : Color from Draw)
    returns mutable DrawableC2D from TestTopOpeDraw;

    Create (C : Curve from Geom2d; CColor : Color from Draw;
    	    Text : CString; TextColor : Color from Draw)
    returns mutable DrawableC2D from TestTopOpeDraw;

    Create (C : Curve from Geom2d; CColor : Color from Draw;
    	    Text : CString; TextColor : Color from Draw;
    	    Discret : Integer;
    	    DispOrigin : Boolean = Standard_True;
            DispCurvRadius : Boolean = Standard_False;
	    RadiusMax : Real = 1.0e3;
	    RatioOfRadius : Real = 0.1)
    returns mutable DrawableC2D from TestTopOpeDraw;

    Pnt2d(me) returns Pnt2d from gp is virtual;
    
    ChangePnt2d(me : mutable; P : Pnt2d);
    
    ChangeCurve(me : mutable; C : Curve from Geom2d);
    
    ChangeText(me : mutable; T : CString from Standard);
    
    Name(me : mutable; N : CString) is redefined;
    
    Whatis(me; I : in out Interpretor from Draw) is redefined;
    ---Purpose: For variable whatis command.

    DrawOn(me; dis : in out Display from Draw) is redefined;
    
fields

    myText2D : Text2D from Draw is protected;
    myText : CString from Standard is protected;
    myTextColor : Color from Draw;

end DrawableC2D;
