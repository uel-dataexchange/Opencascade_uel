-- File:        CurveStyleFont.cdl
-- Created:     Mon Dec  4 12:02:25 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWCurveStyleFont from RWStepVisual

	---Purpose : Read & Write Module for CurveStyleFont

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     CurveStyleFont from StepVisual,
     EntityIterator from Interface

is

	Create returns RWCurveStyleFont;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable CurveStyleFont from StepVisual);

	WriteStep (me; SW : in out StepWriter; ent : CurveStyleFont from StepVisual);

	Share(me; ent : CurveStyleFont from StepVisual; iter : in out EntityIterator);

end RWCurveStyleFont;
