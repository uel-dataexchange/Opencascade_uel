-- File:	ToolPolygon.cdl
-- Created:	Fri Aug  2 08:18:37 1991
-- Author:	Didier PIFFAULT
--		<dpf@sdsun2>
---Copyright:	 Matra Datavision 1991, 1992


generic class ToolPolygon from Intf 
    	    (Point as any;        --  as Pnt2d, Pnt from gp
    	     Polygon as any;
    	     BoundingBox as any)  --  as Box2d, Box from Bnd

	---Purpose: Describes the necessary information about a polyline to
	--          compute the interference between two polylines.

raises  OutOfRange from Standard


is  Bounding       (myclass; thePolyg : Polygon)
    	    	    returns BoundingBox;
    ---Purpose: Returns the bounding box of the polygon.

    DeflectionOverEstimation
		   (myclass; thePolyg : Polygon)
    	    	    returns Real from Standard;
    ---Purpose: Returns the tolerance of the polygon.

    Closed         (myclass; thePolyg : Polygon)
    	    	    returns Boolean from Standard;
    ---Purpose: Returns True if the polyline is closed.

    NbSegments     (myclass; thePolyg : Polygon)
    	    	    returns Integer;
    ---Purpose: Returns the number of Segments in the polyline.
    
    BeginOfSeg     (myclass; thePolyg : Polygon;
    	    	    Index : in Integer)
    	    	    returns Point
    	    	    raises OutOfRange from Standard;
    ---Purpose: Returns the first point of segment of range  <Index> in the
    --          Polygon.

    EndOfSeg       (myclass; thePolyg : Polygon;
    	    	    Index : in Integer)
    	    	    returns Point
    	    	    raises OutOfRange from Standard;
    ---Purpose: Returns the Second point  of the segment  of range Index in
    --          the Polygon.
		 
end ToolPolygon;
