-- File:        ApplicationContext.cdl
-- Created:     Mon Dec  4 12:02:23 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWApplicationContext from RWStepBasic

	---Purpose : Read & Write Module for ApplicationContext

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     ApplicationContext from StepBasic

is

	Create returns RWApplicationContext;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable ApplicationContext from StepBasic);

	WriteStep (me; SW : in out StepWriter; ent : ApplicationContext from StepBasic);

end RWApplicationContext;
