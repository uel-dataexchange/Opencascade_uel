-- File:	TShell.cdl
-- Created:	Mon Dec 17 11:18:44 1990
-- Author:	Remi Lequette
--		<rle@topsn3>
---Copyright:	 Matra Datavision 1990, 1992



class TShell from PTopoDS inherits TShape from PTopoDS

	---Purpose: A topological  Shell shape.

uses
    ShapeEnum from TopAbs

is
    Create returns mutable TShell from PTopoDS;
    	---Level: Internal 
    	
    ShapeType(me) returns ShapeEnum from TopAbs;
    	---Level: Internal 

end TShell;
