-- File:        CsgSolid.cdl
-- Created:     Mon Dec  4 12:02:25 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWCsgSolid from RWStepShape

	---Purpose : Read & Write Module for CsgSolid

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     CsgSolid from StepShape,
     EntityIterator from Interface

is

	Create returns RWCsgSolid;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable CsgSolid from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : CsgSolid from StepShape);

	Share(me; ent : CsgSolid from StepShape; iter : in out EntityIterator);

end RWCsgSolid;
